/******************************************************************************************/
/* 240x240 ST7789 mini display project                Ver.2021-06-03a Kise Kenji, ArchLab */
/******************************************************************************************/
`default_nettype none
/******************************************************************************************/
// 50MHz clock signal of SPI

module SegmentPuzzleProblem0(w_clk, sw_state, enable);
    input wire w_clk, enable;
    input wire [15:0]  sw_state;
    reg [7:0] display_state[3:0];
    wire is_completed = display_state[0][6:0] == 7'b0 &
                        display_state[1][6:0] == 7'b0 &
                        display_state[2][6:0] == 7'b0 &
                        display_state[3][6:0] == 7'b0;

    reg [15:0] timelimit = 60;

    // 0: on
    // 1: off
    always @(posedge w_clk) if(enable) begin
        display_state[0][0] <= ~(0 ^ sw_state[0] ^ sw_state[7] ^ sw_state[14]);
        display_state[0][1] <= ~(0 ^ sw_state[1] ^ sw_state[8] ^ sw_state[15]);
        display_state[0][2] <= ~(0 ^ sw_state[2] ^ sw_state[9]);
        display_state[0][3] <= ~(0 ^ sw_state[3] ^ sw_state[10]);
        display_state[0][4] <= ~(0 ^ sw_state[4] ^ sw_state[11]);
        display_state[0][5] <= ~(0 ^ sw_state[5] ^ sw_state[12]);
        display_state[0][6] <= ~(0 ^ sw_state[6] ^ sw_state[13]);
        display_state[1][0] <= 0;
        display_state[1][1] <= 0;
        display_state[1][2] <= 0;
        display_state[1][3] <= 0;
        display_state[1][4] <= 0;
        display_state[1][5] <= 0;
        display_state[1][6] <= 0;
        display_state[2][0] <= 0;
        display_state[2][1] <= 0;
        display_state[2][2] <= 0;
        display_state[2][3] <= 0;
        display_state[2][4] <= 0;
        display_state[2][5] <= 0;
        display_state[2][6] <= 0;
        display_state[3][0] <= 0;
        display_state[3][1] <= 0;
        display_state[3][2] <= 0;
        display_state[3][3] <= 0;
        display_state[3][4] <= 0;
        display_state[3][5] <= 0;
        display_state[3][6] <= 0;

        display_state[0][7] <= 1;
        display_state[1][7] <= 1;
        display_state[2][7] <= 1;
        display_state[3][7] <= 1;
    end
endmodule

module SegmentPuzzleProblem1(w_clk, sw_state, enable);
    input wire w_clk, enable;
    input wire [15:0]  sw_state;
    reg [7:0] display_state[3:0];
    wire is_completed = display_state[0][6:0] == 7'b0 &
                        display_state[1][6:0] == 7'b0 &
                        display_state[2][6:0] == 7'b0 &
                        display_state[3][6:0] == 7'b0;

    reg [15:0] timelimit = 120;

    // 0: on
    // 1: off
    always @(posedge w_clk) if(enable) begin
        display_state[0][0] <= ~(0 ^ sw_state[0] ^ sw_state[11] ^ sw_state[13]);
        display_state[0][1] <= ~(0 ^ sw_state[3] ^ sw_state[7]);
        display_state[0][2] <= ~(0 ^ sw_state[4] ^ sw_state[9]);
        display_state[0][3] <= ~(0 ^ sw_state[2] ^ sw_state[12] ^ sw_state[15]);
        display_state[0][4] <= ~(0 ^ sw_state[6] ^ sw_state[10]);
        display_state[0][5] <= ~(0 ^ sw_state[5] ^ sw_state[8]);
        display_state[0][6] <= ~(0 ^ sw_state[1] ^ sw_state[14]);
        display_state[1][0] <= ~(0 ^ sw_state[0] ^ sw_state[12]);
        display_state[1][1] <= ~(0 ^ sw_state[3] ^ sw_state[8]);
        display_state[1][2] <= ~(0 ^ sw_state[4] ^ sw_state[10]);
        display_state[1][3] <= ~(0 ^ sw_state[2] ^ sw_state[11] ^ sw_state[14]);
        display_state[1][4] <= ~(0 ^ sw_state[6] ^ sw_state[9]);
        display_state[1][5] <= ~(0 ^ sw_state[5] ^ sw_state[7]);
        display_state[1][6] <= ~(0 ^ sw_state[1] ^ sw_state[13] ^ sw_state[15]);
        display_state[2][0] <= 0;
        display_state[2][1] <= 0;
        display_state[2][2] <= 0;
        display_state[2][3] <= 0;
        display_state[2][4] <= 0;
        display_state[2][5] <= 0;
        display_state[2][6] <= 0;
        display_state[3][0] <= 0;
        display_state[3][1] <= 0;
        display_state[3][2] <= 0;
        display_state[3][3] <= 0;
        display_state[3][4] <= 0;
        display_state[3][5] <= 0;
        display_state[3][6] <= 0;

        display_state[0][7] <= 1;
        display_state[1][7] <= 1;
        display_state[2][7] <= 1;
        display_state[3][7] <= 1;
   end
endmodule

module SegmentPuzzleProblem2(w_clk, sw_state, enable);
    input wire w_clk, enable;
    input wire [15:0]  sw_state;
    reg [7:0] display_state[3:0];
    wire is_completed = display_state[0][6:0] == 7'b0 &
                        display_state[1][6:0] == 7'b0 &
                        display_state[2][6:0] == 7'b0 &
                        display_state[3][6:0] == 7'b0;

    reg [15:0] timelimit = 180;

    // 0: on
    // 1: off
    always @(posedge w_clk) if(enable) begin
        display_state[0][0] <= ~(0 ^ sw_state[14]);
        display_state[0][1] <= ~(0 ^ sw_state[0] ^ sw_state[3] ^ sw_state[9] ^ sw_state[11]);
        display_state[0][2] <= ~(0 ^ sw_state[0] ^ sw_state[1] ^ sw_state[9]);
        display_state[0][3] <= ~(0 ^ sw_state[4] ^ sw_state[14] ^ sw_state[15]);
        display_state[0][4] <= ~(0 ^ sw_state[3] ^ sw_state[5] ^ sw_state[6] ^ sw_state[14]);
        display_state[0][5] <= ~(0 ^ sw_state[6] ^ sw_state[8] ^ sw_state[13] ^ sw_state[14]);
        display_state[0][6] <= ~(0 ^ sw_state[0]);
        display_state[1][0] <= ~(0 ^ sw_state[0] ^ sw_state[11] ^ sw_state[12]);
        display_state[1][1] <= ~(0 ^ sw_state[2] ^ sw_state[6]);
        display_state[1][2] <= ~(0 ^ sw_state[1] ^ sw_state[2] ^ sw_state[3] ^ sw_state[5] ^ sw_state[9]);
        display_state[1][3] <= ~(0 ^ sw_state[0] ^ sw_state[6] ^ sw_state[8]);
        display_state[1][4] <= ~(0 ^ sw_state[2] ^ sw_state[3]);
        display_state[1][5] <= ~(0 ^ sw_state[2] ^ sw_state[7] ^ sw_state[9] ^ sw_state[11]);
        display_state[1][6] <= ~(0 ^ sw_state[2]);
        display_state[2][0] <= ~(0 ^ sw_state[2] ^ sw_state[3] ^ sw_state[11] ^ sw_state[12]);
        display_state[2][1] <= ~(0 ^ sw_state[4] ^ sw_state[6] ^ sw_state[6] ^ sw_state[8] ^ sw_state[10] ^ sw_state[14]);
        display_state[2][2] <= ~(0 ^ sw_state[3] ^ sw_state[5] ^ sw_state[9] ^ sw_state[14]);
        display_state[2][3] <= ~(0 ^ sw_state[2] ^ sw_state[15]);
        display_state[2][4] <= ~(0 ^ sw_state[9] ^ sw_state[14]);
        display_state[2][5] <= ~(0 ^ sw_state[14]);
        display_state[2][6] <= ~(0 ^ sw_state[2] ^ sw_state[7]);
        display_state[3][0] <= 0;
        display_state[3][1] <= 0;
        display_state[3][2] <= 0;
        display_state[3][3] <= 0;
        display_state[3][4] <= 0;
        display_state[3][5] <= 0;
        display_state[3][6] <= 0;

        display_state[0][7] <= 1;
        display_state[1][7] <= 1;
        display_state[2][7] <= 1;
        display_state[3][7] <= 1;
   end
endmodule


module SegmentPuzzleProblem3(w_clk, sw_state, enable);
    input wire w_clk, enable;
    input wire [15:0]  sw_state;
    reg [7:0] display_state[3:0];
    wire is_completed = display_state[0][6:0] == 7'b0 &
                        display_state[1][6:0] == 7'b0 &
                        display_state[2][6:0] == 7'b0 &
                        display_state[3][6:0] == 7'b0;

    reg [15:0] timelimit = 900;

    // 0: on
    // 1: off
    always @(posedge w_clk) if(enable) begin
        display_state[0][0] <= ~(0 ^ sw_state[2] ^ sw_state[6] ^ sw_state[7] ^ sw_state[14]);
        display_state[0][1] <= ~(0 ^ sw_state[0] ^ sw_state[4] ^ sw_state[7] ^ sw_state[11] ^ sw_state[12] ^ sw_state[13]);
        display_state[0][2] <= ~(0 ^ sw_state[6] ^ sw_state[8] ^ sw_state[9] ^ sw_state[11]);
        display_state[0][3] <= ~(0 ^ sw_state[1] ^ sw_state[11] ^ sw_state[12]);
        display_state[0][4] <= ~(0 ^ sw_state[3] ^ sw_state[12] ^ sw_state[15]);
        display_state[0][5] <= ~(0 ^ sw_state[4] ^ sw_state[5] ^ sw_state[6] ^ sw_state[7] ^ sw_state[8] ^ sw_state[9] ^ sw_state[10] ^ sw_state[14]);
        display_state[0][6] <= ~(0 ^ sw_state[0] ^ sw_state[1]);
        display_state[1][0] <= ~(0 ^ sw_state[3] ^ sw_state[15]);
        display_state[1][1] <= ~(0 ^ sw_state[3] ^ sw_state[4] ^ sw_state[14]);
        display_state[1][2] <= ~(0 ^ sw_state[1] ^ sw_state[4] ^ sw_state[5] ^ sw_state[9] ^ sw_state[10] ^ sw_state[12]);
        display_state[1][3] <= ~(0 ^ sw_state[6] ^ sw_state[8] ^ sw_state[11] ^ sw_state[15]);
        display_state[1][4] <= ~(0 ^ sw_state[2] ^ sw_state[5] ^ sw_state[7] ^ sw_state[8] ^ sw_state[10] ^ sw_state[13]);
        display_state[1][5] <= ~(0 ^ sw_state[4] ^ sw_state[9]);
        display_state[1][6] <= ~(0 ^ sw_state[0] ^ sw_state[8] ^ sw_state[14]);
        display_state[2][0] <= ~(0 ^ sw_state[1] ^ sw_state[2] ^ sw_state[4] ^ sw_state[6]);
        display_state[2][1] <= ~(0 ^ sw_state[0] ^ sw_state[10] ^ sw_state[11] ^ sw_state[13]);
        display_state[2][2] <= ~(0 ^ sw_state[0] ^ sw_state[2] ^ sw_state[5] ^ sw_state[8] ^ sw_state[12]);
        display_state[2][3] <= ~(0 ^ sw_state[3]);
        display_state[2][4] <= ~(0 ^ sw_state[1] ^ sw_state[7] ^ sw_state[13]);
        display_state[2][5] <= ~(0 ^ sw_state[10] ^ sw_state[14] ^ sw_state[15]);
        display_state[2][6] <= ~(0 ^ sw_state[5] ^ sw_state[9]);
        display_state[3][0] <= ~(0 ^ sw_state[1] ^ sw_state[4] ^ sw_state[5] ^ sw_state[6] ^ sw_state[7] ^ sw_state[8] ^ sw_state[13] ^ sw_state[14] ^ sw_state[15]);
        display_state[3][1] <= ~(0 ^ sw_state[2] ^ sw_state[3]);
        display_state[3][2] <= ~(0 ^ sw_state[6] ^ sw_state[11] ^ sw_state[12] ^ sw_state[15]);
        display_state[3][3] <= ~(0 ^ sw_state[6] ^ sw_state[9] ^ sw_state[10] ^ sw_state[12]);
        display_state[3][4] <= ~(0 ^ sw_state[4] ^ sw_state[12]);
        display_state[3][5] <= ~(0 ^ sw_state[3] ^ sw_state[8]);
        display_state[3][6] <= ~(0 ^ sw_state[0] ^ sw_state[5] ^ sw_state[10]);

        display_state[0][7] <= 1;
        display_state[1][7] <= 1;
        display_state[2][7] <= 1;
        display_state[3][7] <= 1;
    end
endmodule


module SecCounter(w_clk, enable, reset);
    input wire w_clk, enable, reset;

    reg[31:0] clk_count = 0;
    reg[31:0] elapsed_sec = 0;
    always @(posedge w_clk) begin
        clk_count   <= reset ? 0 : (~enable) ? clk_count   : (clk_count+1 == 100_000_000 ? 0 : clk_count + 1);
        elapsed_sec <= reset ? 0 : (~enable) ? elapsed_sec : (clk_count+1 == 100_000_000 ? elapsed_sec+1 : elapsed_sec);
    end
endmodule

module Timer(preset_time_sec, w_clk, enable, reset);
    input wire[15:0] preset_time_sec;
    input wire w_clk, enable, reset;

    SecCounter counter(w_clk, enable, reset);

    reg [15:0] remaining_time_sec;
    reg is_finished;

    always @(posedge w_clk) begin
        remaining_time_sec <= reset ? preset_time_sec : (preset_time_sec > counter.elapsed_sec ? preset_time_sec - counter.elapsed_sec : 0);
        is_finished <= remaining_time_sec == 0;
    end
endmodule

function [7:0] ConvertDigitTo7SegDisplayState;
    input [3:0] digit;

    case (digit)
        4'd0: ConvertDigitTo7SegDisplayState = 8'b11000000;  // 0
        4'd1: ConvertDigitTo7SegDisplayState = 8'b11111001;  // 1
        4'd2: ConvertDigitTo7SegDisplayState = 8'b10100100;  // 2
        4'd3: ConvertDigitTo7SegDisplayState = 8'b10110000;  // 3
        4'd4: ConvertDigitTo7SegDisplayState = 8'b10011001;  // 4
        4'd5: ConvertDigitTo7SegDisplayState = 8'b10010010;  // 5
        4'd6: ConvertDigitTo7SegDisplayState = 8'b10000010;  // 6
        4'd7: ConvertDigitTo7SegDisplayState = 8'b11111000;  // 7
        4'd8: ConvertDigitTo7SegDisplayState = 8'b10000000;  // 8
        4'd9: ConvertDigitTo7SegDisplayState = 8'b10010000;  // 9
        default: ConvertDigitTo7SegDisplayState = 8'b11111111; // すべてオフ（エラーケース）
    endcase
endfunction

module TimeTo7SegDisplayStateConverter(w_clk, time_sec);
    input wire w_clk;
    input wire[15:0] time_sec;

    reg [3:0] digits[3:0];
    wire [7:0] display_state[3:0];

    always @(posedge w_clk) begin
        digits[0] = time_sec % 10;
        digits[1] = (time_sec / 10) % 6;
        digits[2] = (time_sec / 60) % 10;
        digits[3] = (time_sec / 600) % 6;
    end
    assign display_state[0] = ConvertDigitTo7SegDisplayState(digits[0]);
    assign display_state[1] = ConvertDigitTo7SegDisplayState(digits[1]);
    assign display_state[2] = ConvertDigitTo7SegDisplayState(digits[2]);
    assign display_state[3] = ConvertDigitTo7SegDisplayState(digits[3]);

endmodule

module GameState(
        w_clk,
        sw,
        is_pressed_left_btn,
        is_pressed_right_btn,
        is_pressed_top_btn,
        is_pressed_bottom_btn,
        is_pressed_center_btn
);
    input  wire w_clk;
    input  wire is_pressed_left_btn, is_pressed_right_btn, is_pressed_top_btn, is_pressed_bottom_btn, is_pressed_center_btn;

    input  wire [15:0]  sw;

    SegmentPuzzleProblem0 problem0(w_clk, sw, (~game_finished));
    SegmentPuzzleProblem1 problem1(w_clk, sw, (~game_finished));
    SegmentPuzzleProblem2 problem2(w_clk, sw, (~game_finished));
    SegmentPuzzleProblem3 problem3(w_clk, sw, (~game_finished));

    wire problem_completed = game_mode == 0 ? problem0.is_completed :
                             game_mode == 1 ? problem1.is_completed :
                             game_mode == 2 ? problem2.is_completed :
                             game_mode == 3 ? problem3.is_completed :
                                              0;

    reg game_finished = 0;
    reg game_started = 0;
    reg reset_game = 0;
    reg[1:0] game_mode = 0;
    always @(posedge w_clk) begin
        game_mode = game_started ? game_mode :
                    is_pressed_top_btn    ? 0 :
                    is_pressed_left_btn   ? 1 :
                    is_pressed_center_btn ? 2 :
                    is_pressed_right_btn  ? 3 :
                    game_mode;
        reset_game = is_pressed_bottom_btn;
        game_started = (~reset_game) & (game_started | is_pressed_top_btn | is_pressed_left_btn | is_pressed_center_btn | is_pressed_right_btn);
        game_finished = game_started & (game_finished | problem_completed | timer.is_finished);

    end

    wire [15:0] timelimit = game_mode == 0 ? problem0.timelimit :
                            game_mode == 1 ? problem1.timelimit :
                            game_mode == 2 ? problem2.timelimit :
                            game_mode == 3 ? problem3.timelimit :
                                             0;

    Timer timer(timelimit, w_clk, game_started & (~game_finished), reset_game);
    TimeTo7SegDisplayStateConverter converter(w_clk, timer.remaining_time_sec);

    // controll display
    reg[31:0] clk_count = 0;
    always @(posedge w_clk) begin
        clk_count <= (clk_count == 1_600_000 ? 0 : clk_count + 1);
    end

    wire [2:0] target_seg_display_idx = (clk_count / 200_000);
    wire [7:0] is_lighted_seg_display = ~(1<<target_seg_display_idx);
    wire [7:0] seg_display_state = (~game_started) ? 0 :
                                   target_seg_display_idx >= 4 ? converter.display_state[target_seg_display_idx-4] :
                                   game_mode == 0 ? problem0.display_state[target_seg_display_idx] :
                                   game_mode == 1 ? problem1.display_state[target_seg_display_idx] :
                                   game_mode == 2 ? problem2.display_state[target_seg_display_idx] :
                                   game_mode == 3 ? problem3.display_state[target_seg_display_idx] :
                                                    0;
endmodule

/******************************************************************************************/
module m_main(
        w_clk,
        st7789_SDA,
        st7789_SCL,
        st7789_DC,
        st7789_RES,
        led,
        sw,
        is_pressed_left_btn,
        is_pressed_right_btn,
        is_pressed_top_btn,
        is_pressed_bottom_btn,
        is_pressed_center_btn,
        seg_display_state,
        is_lighted_seg_display
);
    input  wire w_clk; // main clock signal (100MHz)
    output wire st7789_SCL;
    inout  wire st7789_SDA;
    output wire st7789_DC;
    output wire st7789_RES;
    output wire [15:0] led;
    input  wire [15:0] sw;
    input  wire is_pressed_left_btn, is_pressed_right_btn, is_pressed_top_btn, is_pressed_bottom_btn, is_pressed_center_btn;
    output wire [7:0] seg_display_state;
    output wire [7:0] is_lighted_seg_display;

    GameState game_state(
            w_clk,
            sw,
            is_pressed_left_btn,
            is_pressed_right_btn,
            is_pressed_top_btn,
            is_pressed_bottom_btn,
            is_pressed_center_btn
    );
    assign seg_display_state = game_state.seg_display_state;
    assign is_lighted_seg_display = game_state.is_lighted_seg_display;


    wire w_clk_t = w_clk;
    reg [15:0] r_sw=0;
    always @(posedge w_clk_t) r_sw <= sw;
    /**********************************************************************************/
    reg [7:0] r_x=0, r_y=0;
    always @(posedge w_clk_t) begin
        r_x <= (r_x==239) ? 0 : r_x + 1;
        r_y <= (r_y==239) ? 0 : (r_x==239) ? r_y + 1 : r_y;
    end

    reg [15:0] r_st_wadr  = 0; //{ r_y[7:0], r_sx[7:0]};
    reg        r_st_we    = 0; // cam_we && (r_sx<256) && (r_y<256);
    reg [15:0] r_st_wdata = 0; // cam_dout;
    always @(posedge w_clk_t) r_st_wadr  <= {r_y, r_x};
    always @(posedge w_clk_t) r_st_we    <= 1;

    always @(posedge w_clk_t) r_st_wdata <= game_state.game_finished ? (game_state.problem_completed ? image_succeeded[r_st_wadr] : image_failed[r_st_wadr]) :
                                            game_state.game_started  ? image_start[r_st_wadr] :
                                                                       image_start[r_st_wadr];

    reg [15:0] vmem [0:65535]; // video memory, 256 x 256 (65,536) x 12bit color
    always @(posedge w_clk_t) if(r_st_we) vmem[r_st_wadr] <= r_st_wdata;

    wire [15:0] w_raddr;
    reg [15:0] r_rdata = 0;
    reg [15:0] r_raddr = 0;
    always @(posedge w_clk_t) r_raddr <= w_raddr;
    always @(posedge w_clk_t) r_rdata <= vmem[r_raddr];

    wire [1:0] w_mode = 2'b11;
    m_st7789_display display0 (w_clk_t, st7789_SDA, st7789_SCL, st7789_DC, st7789_RES, w_raddr, r_rdata, w_mode);

    reg [15:0] image_start [0:65535] = {
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hF71C, 16'hD618, 16'hD658, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hF79D, 16'hF71C, 16'hD5D7, 16'hBC93, 16'hC4D3, 16'hC492, 16'hA30D, 16'hAB8E, 16'hE618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'hD5D8, 16'hB451, 16'hB3CF, 16'hB3CF, 16'hCCD3, 16'hC451, 16'hAB8E, 16'h9B0C, 16'hBC10, 16'hC493, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hE6DB, 16'hD618, 16'hB492, 16'hA34D, 16'hBC52, 16'hCCD4, 16'hDD97, 16'hEE18, 16'hC493, 16'h8A8A, 16'h928A, 16'h928A, 16'h8A89, 16'hB3CF, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hF71C, 16'hD5D7, 16'hBC92, 16'hA38F, 16'hB411, 16'hCCD5, 16'hDD97, 16'hEE19, 16'hEE19, 16'hE5D8, 16'hB410, 16'h79C6, 16'hBC10, 16'hC451, 16'hBC10, 16'h9B0C, 16'hAB4D, 16'hEE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hEEDB, 16'hDDD8, 16'hC493, 16'hC493, 16'hC493, 16'hD515, 16'hE5D8, 16'hE5D9, 16'hEE1A, 16'hE61A, 16'hE619, 16'hEDD8, 16'hABCF, 16'h81C6, 16'hBC10, 16'hDD56, 16'hDD15, 16'hC410, 16'hAB4D, 16'hB38E, 16'hE659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hE69A, 16'hD597, 16'hB411, 16'hBC52, 16'hCCD4, 16'hDD57, 16'hDD98, 16'hEE19, 16'hEE1A, 16'hE619, 16'hE619, 16'hE5D9, 16'hE619, 16'hE5D8, 16'hA38E, 16'h8A49, 16'hD4D3, 16'hDD56, 16'hDD56, 16'hDD55, 16'hCCD3, 16'hDD14, 16'hC410, 16'hD596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hE659, 16'hD556, 16'hB410, 16'hAB8F, 16'hCC93, 16'hD515, 16'hE598, 16'hE619, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE598, 16'hA34D, 16'h8A49, 16'hD514, 16'hDD96, 16'hDD56, 16'hDD56, 16'hDD55, 16'hDD55, 16'hE596, 16'hC451, 16'hC4D4, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hCD55, 16'hC492, 16'hA34E, 16'hBC11, 16'hC493, 16'hDD97, 16'hE5D9, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE619, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE619, 16'hE619, 16'hE5D8, 16'hA34E, 16'h8A89, 16'hD514, 16'hDD96, 16'hDD55, 16'hDD55, 16'hDD56, 16'hDD56, 16'hDD56, 16'hDD96,
        16'hC451, 16'hBC51, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hDE18, 16'hC4D4, 16'hA2CC, 16'hAB4D, 16'hCCD4, 16'hDD97, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hE61A, 16'hE619, 16'hE619, 16'hE619, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hEDD8, 16'hAB8F, 16'h8A8A, 16'hCCD3, 16'hDD96, 16'hDD55, 16'hDD96, 16'hDD56, 16'hDD56, 16'hDD56, 16'hDD56, 16'hDD96, 16'hCCD3, 16'hB3D0, 16'hFF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hC514, 16'hA34D, 16'hAB0D, 16'hBC51, 16'hDD56, 16'hEE19, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE619, 16'hE61A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hEDD8,
        16'hA38E, 16'h8A49, 16'hD514, 16'hDD96, 16'hD556, 16'hDD96, 16'hDD96, 16'hDD56, 16'hDD56, 16'hDD56, 16'hDD96, 16'hDD96, 16'hDD55, 16'hAB8E, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD618, 16'hB492, 16'h9ACB, 16'hB34E, 16'hD4D4, 16'hE598, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE619, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE61A, 16'hEE1A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hEE19, 16'hABCF, 16'h8249, 16'hCCD3, 16'hDD96, 16'hD556, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD56, 16'hDD56, 16'hDD56, 16'hDD96, 16'hDD96, 16'hDD96, 16'hAB4D, 16'hE65A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75C, 16'hCD96, 16'h9B4C, 16'h92CB, 16'hC492, 16'hD556, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hEE1A, 16'hEE1A,
        16'hEE1A, 16'hEE19, 16'hEE19, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hBC52, 16'h8A49, 16'hCCD3, 16'hDD96, 16'hD555, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD56, 16'hDD56, 16'hDD96, 16'hDD96, 16'hDD96, 16'hE597, 16'hAB8E, 16'hDE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DA, 16'hB4D2, 16'h8208, 16'hAB8E, 16'hC4D3, 16'hE619, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE619, 16'hEE1A, 16'hC494, 16'h81C8, 16'hCC92, 16'hDD96, 16'hDD56, 16'hDD56, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD56, 16'hDD56, 16'hDD96, 16'hDD96, 16'hDD96, 16'hE5D7, 16'hB3CF, 16'hD5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hB451, 16'h8A49, 16'hB3D0, 16'hCD15, 16'hE619,
        16'hEE5A, 16'hEE1A, 16'hE619, 16'hE619, 16'hEE19, 16'hEE1A, 16'hEE19, 16'hE619, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE619, 16'hEE1A, 16'hD556, 16'h9249, 16'hC452, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hE5D7, 16'hB3D0, 16'hCD56, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hDE18, 16'hB451, 16'h8A09, 16'hA34E, 16'hD556, 16'hEE1A, 16'hEE5A, 16'hEE1A, 16'hE619, 16'hE619, 16'hE61A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hE61A, 16'hE61A, 16'hE619, 16'hEE5A, 16'hD556, 16'h928B, 16'hBC11, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hE5D7, 16'hBC11, 16'hC555, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hDE59, 16'hA3CE, 16'h7905, 16'hAB8F, 16'hDD57, 16'hEE19, 16'hEE5A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE619, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hE61A, 16'hE619, 16'hEE1A, 16'hDD97, 16'hA34E, 16'hAB8E, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD56, 16'hDD56, 16'hDD96, 16'hDD96, 16'hDD96, 16'hE5D7, 16'hBC11, 16'hC514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hA410, 16'h8A08, 16'hB3D1, 16'hDD97, 16'hE619, 16'hEE5A, 16'hE619, 16'hEE19, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE619, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hE619, 16'hEE5A, 16'hDD97, 16'h9B0C, 16'hA34D, 16'hDD56, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD56,
        16'hDD56, 16'hDD96, 16'hDD96, 16'hDD96, 16'hE5D7, 16'hBC51, 16'hBCD4, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hB492, 16'h924A, 16'hB3D1, 16'hD557, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE619, 16'hE619, 16'hEE1A, 16'hEE1A, 16'hE61A, 16'hE619, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hE619, 16'hE61A, 16'hE5D8, 16'hAB8F, 16'h92CB, 16'hDD55, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hE5D7, 16'hC451, 16'hC514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hC595, 16'h9B0B, 16'hAB8E, 16'hD556, 16'hEE19, 16'hEE1A, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hE619, 16'hE619, 16'hEE19, 16'hB3D0, 16'h9ACC, 16'hDD15, 16'hDD96,
        16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD56, 16'hDD96, 16'hDD96, 16'hDD96, 16'hE5D7, 16'hC492, 16'hBCD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hCD55, 16'hA34D, 16'hAB8E, 16'hCD15, 16'hE5D9, 16'hEE1A, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hE619, 16'hE619, 16'hEE1A, 16'hBC52, 16'h9249, 16'hCCD3, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD56, 16'hDD56, 16'hDD96, 16'hDD96, 16'hDD97, 16'hE5D7, 16'hBC11, 16'hBCD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD5D7, 16'hB38E, 16'hAB0D, 16'hCC94, 16'hE5D9, 16'hEE1A, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hEE1A,
        16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hE619, 16'hEE1A, 16'hCC93, 16'h928A, 16'hC492, 16'hE596, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD56, 16'hDD56, 16'hDD96, 16'hDD96, 16'hDD96, 16'hE5D7, 16'hC452, 16'hC555, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'hB3CF, 16'hA2CB, 16'hC452, 16'hE5D8, 16'hEE1A, 16'hE61A, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hE619, 16'hEE5A, 16'hD515, 16'h8A49, 16'hBC11, 16'hE597, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD56, 16'hDD56, 16'hDD96, 16'hDD96, 16'hDD97, 16'hE5D7, 16'hC452, 16'hCD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hC4D3, 16'h9A49, 16'hB38F, 16'hDD56, 16'hEE1A, 16'hE61A, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619,
        16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hE61A, 16'hE619, 16'hEE5A, 16'hD515, 16'h8A49, 16'hBC52, 16'hE5D7, 16'hE5D7, 16'hDD97, 16'hDDD6, 16'hDDD6, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD56, 16'hDD56, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD97, 16'hE5D7, 16'hBC10, 16'hCD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hC596, 16'h92CB, 16'h9A8B, 16'hD4D4, 16'hEE19, 16'hEE1A, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE619, 16'hD516, 16'hA30C, 16'hCCD3, 16'hEE18, 16'hDD56, 16'hDD55, 16'hDD56, 16'hDD55, 16'hD514, 16'hDD55, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD56, 16'hDD56, 16'hDD96, 16'hDD96, 16'hDD56, 16'hDD56, 16'hDD56, 16'hDD96, 16'hDD96, 16'hDD97, 16'hDD97, 16'hE5D7, 16'hBC11, 16'hDDD7, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9A, 16'hA38E, 16'h9249, 16'hCC93, 16'hE598, 16'hEE1A, 16'hE619, 16'hE619, 16'hE619, 16'hE619,
        16'hE61A, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hEE1A, 16'hDD97, 16'h7986, 16'h8A08, 16'hB38E, 16'hB3CF, 16'hC451, 16'hBBD0, 16'hB38E, 16'hB38E, 16'hA30C, 16'hAB8E, 16'hBC10, 16'hCCD4, 16'hDD96, 16'hDD56, 16'hDD56, 16'hDD56, 16'hDD56, 16'hDD96, 16'hDD56, 16'hDD56, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD97, 16'hDD97, 16'hE5D7, 16'hBC10, 16'hDE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD96, 16'h9248, 16'hB34E, 16'hDD16, 16'hEE1A, 16'hE61A, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hEE5A, 16'hCD15, 16'h8249, 16'hC514, 16'hE69A, 16'hF75D, 16'hFF5E, 16'hFF5E, 16'hE65A, 16'hDD55, 16'hDD96, 16'hDD55, 16'hD515, 16'hDD55, 16'hDD96, 16'hDD56, 16'hDD56, 16'hDD56, 16'hDD56,
        16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD97, 16'hDD97, 16'hDD97, 16'hE5D7, 16'hB410, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF79E, 16'hEF1C, 16'hEF1C, 16'hEEDC, 16'hE65A, 16'hDE19, 16'hDE19, 16'hD5D8, 16'hCD96, 16'hDE18, 16'hD5D8, 16'hD5D7, 16'hDE59, 16'hE659, 16'hE65A, 16'hEEDC, 16'hF71C, 16'hF75D, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB,
        16'hAC10, 16'h8A08, 16'hCC93, 16'hEDD8, 16'hEE19, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE61A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE61A, 16'hE5D9, 16'hD515, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF6DB, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD56, 16'hDD56, 16'hDD56, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD97, 16'hDD97, 16'hE597, 16'hE597, 16'hDD97, 16'hB3D0, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hEF1C, 16'hDE59, 16'hD596, 16'hB451, 16'hABCF, 16'hABCF, 16'hB38F, 16'hAB4E, 16'hBC10, 16'hB410, 16'hC451, 16'hAB8F, 16'hC493, 16'hB410, 16'hC493, 16'hBC52, 16'hABD0, 16'hB411, 16'hB3D0, 16'hAB8F, 16'h8A8A, 16'hA34D, 16'h9B0D, 16'h934D, 16'hC4D3, 16'hCD14, 16'hDE18, 16'hD5D7, 16'h8A8A, 16'hA2CC, 16'hDD16, 16'hEDD9, 16'hE61A, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE61A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hEE19, 16'hC4D3, 16'hB451, 16'hF6DB, 16'hFF9E, 16'hFFDF, 16'hFFDF,
        16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'hDDD7, 16'hDD56, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDDD7, 16'hDDD7, 16'hE5D7, 16'hDD96, 16'hABCF, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF71C, 16'hDE19, 16'hCD15, 16'hBC11, 16'hB3CF, 16'hAB8E, 16'hA38E, 16'hB410, 16'hCD14, 16'hD596, 16'hDDD8, 16'hDDD8, 16'hE619, 16'hE619, 16'hE5D8, 16'hE619, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDD97, 16'hE5D8, 16'hDDD8,
        16'hE619, 16'hE619, 16'hEE1A, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hBC52, 16'hAB8E, 16'h92CB, 16'h6800, 16'h8145, 16'hBC11, 16'hE598, 16'hEE19, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hEE5A, 16'hCD15, 16'hB411, 16'hEE19, 16'hE618, 16'hEE19, 16'hEE5A, 16'hEE9B, 16'hEE9A, 16'hD597, 16'hEE9B, 16'hF71D, 16'hEE5A, 16'hDD56, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDDD7, 16'hE5D7, 16'hE5D7, 16'hDD96, 16'hB411, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD97, 16'hCD55, 16'hCD55, 16'hD596, 16'hD596, 16'hD596, 16'hD596, 16'hD596, 16'hD5D8, 16'hE659, 16'hE659, 16'hE69A, 16'hEEDB, 16'hEEDB, 16'hEEDC, 16'hF75D, 16'hFF5D, 16'hFF5E, 16'hF75E, 16'hFF5E, 16'hF75D, 16'hFF9E, 16'hFF9E, 16'hF75E, 16'hF75E, 16'hFF9E, 16'hF75E, 16'hFF5E, 16'hFF5E, 16'hF75D, 16'hF75E, 16'hF75D, 16'hFF9E, 16'hFF9F, 16'hFF9E, 16'hFF9F, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hE69A, 16'hCD55, 16'hABCF, 16'hB3CF, 16'hB410, 16'hBC93, 16'hD5D7, 16'hE69A, 16'hF71C, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFF1D, 16'hFEDD, 16'hF69C, 16'hF69B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hEE1A, 16'hE5D9, 16'hE5D8, 16'hDD97, 16'hDD56, 16'hDD15, 16'hCCD4, 16'hCCD4, 16'hE5D8, 16'hF65B, 16'hFE5A, 16'hC452, 16'h824A, 16'h9B0C, 16'hD4D4, 16'hEE19, 16'hEE19, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE1A, 16'hEE1A,
        16'hEE1A, 16'hEE1A, 16'hE619, 16'hEE1A, 16'hE5D8, 16'hA38E, 16'hE5D8, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEDD8, 16'hDD97, 16'hDD56, 16'hDD56, 16'hCCD3, 16'hCCD4, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD96, 16'hDD97, 16'hE5D7, 16'hE5D7, 16'hDDD7, 16'hDDD7, 16'hDDD7, 16'hDDD7, 16'hDDD7, 16'hE5D7, 16'hE5D7, 16'hD555, 16'hB451, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hC493, 16'h924A, 16'h9249, 16'hA30C, 16'hBBD0, 16'hBC11, 16'hB38F, 16'hB34E, 16'hA2CC, 16'hB34E, 16'hAB4D, 16'hAB4D, 16'hB38E, 16'hAB4E, 16'hA30D, 16'hA30D, 16'hAB4E, 16'hA34D, 16'hAB4D, 16'hAB8E, 16'hA30D, 16'hAB8E, 16'hB3D0, 16'hAB8E, 16'hAB8E, 16'hAB8F, 16'hAB8F, 16'hAB8F, 16'hAB4E, 16'h9B0D, 16'hBC11, 16'hA38F, 16'hA38E, 16'hABD0, 16'hABD0, 16'hABD0, 16'hB410, 16'hBC92, 16'hB411, 16'hC4D3, 16'hBC92, 16'hBCD3, 16'hD596, 16'hCD55, 16'hCD96, 16'hD5D7, 16'hDE59, 16'hDE59, 16'hE69A, 16'hEEDB, 16'hEEDB, 16'hF75D, 16'hFF9E, 16'hF79E, 16'hFFDE, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hDE18, 16'hBC92, 16'hA38E, 16'hAB8F, 16'hBC92, 16'hD597, 16'hEEDB, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hF6DC,
        16'hF69B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF69B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hF65A, 16'hF61A, 16'hEDD9, 16'hDD56, 16'hD515, 16'hCCD4, 16'hAB8F, 16'h7985, 16'hABCF, 16'hEDD8, 16'hEE19, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE61A, 16'hEE19, 16'hABD0, 16'hD556, 16'hEE59, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE18, 16'hE5D8, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hDD97, 16'hE597, 16'hE597, 16'hDD96, 16'hDD96, 16'hE596, 16'hE597, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hDDD7, 16'hDDD7, 16'hDDD7, 16'hDDD7, 16'hE5D8, 16'hC4D3, 16'hBC92, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC4D3, 16'hA30D, 16'hAB4E, 16'h9A8A, 16'hB34E, 16'hD515, 16'hEDD9, 16'hE5D8, 16'hE598, 16'hE598, 16'hE598, 16'hE597, 16'hDD97, 16'hE597, 16'hDD56, 16'hD516, 16'hD516, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD514, 16'hD4D4, 16'hD515, 16'hD515, 16'hCCD4, 16'hCCD4, 16'hD514, 16'hD514, 16'hCCD4, 16'hD556, 16'hD555, 16'hCCD4, 16'hC4D4, 16'hCCD3, 16'hC492, 16'hC493, 16'hC492, 16'hBC51, 16'hCC92, 16'hBC51,
        16'hAB8F, 16'hB3CF, 16'hB3CF, 16'hA30D, 16'hA30D, 16'h9B0C, 16'h9ACB, 16'h9ACB, 16'h9B0C, 16'h928A, 16'h9B4C, 16'hA38E, 16'hA38E, 16'hAC10, 16'hC4D3, 16'hBCD3, 16'hC555, 16'hD5D6, 16'hDE18, 16'hE69A, 16'hEF1B, 16'hF75D, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hEEDB, 16'hBC92, 16'h9B0C, 16'h9B4D, 16'hCD56, 16'hE69A, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hF6DC, 16'hF69C, 16'hF69B, 16'hF69B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hEE5A, 16'hF65A, 16'hF61A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hE5D9, 16'hEE1A, 16'hEDD8, 16'hA34E, 16'h8A8B, 16'hDD55, 16'hEE19, 16'hEE1A, 16'hE61A, 16'hE619, 16'hEE1A, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE19, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619,
        16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hEE5A, 16'hC493, 16'hBC52, 16'hEE19, 16'hE618, 16'hE5D8, 16'hEE19, 16'hEE19, 16'hEE19, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D7, 16'hE5D8, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hDDD7, 16'hDDD7, 16'hDDD7, 16'hDDD7, 16'hE618, 16'hBC92, 16'hC514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC555, 16'h924A, 16'hDD15, 16'hDCD4, 16'hC3D1, 16'h9A8B, 16'hC411, 16'hE5D9, 16'hEE1A, 16'hE5D9, 16'hE619, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hE5D9, 16'hE5D9, 16'hE619, 16'hDD97, 16'hD556, 16'hD557, 16'hCD15, 16'hCCD5, 16'hC494, 16'hBC93, 16'hB411, 16'hB3D0, 16'hB3D0, 16'hAB8E, 16'h9B0C, 16'h92CB, 16'h92CB, 16'hA38D, 16'hB450, 16'hAC50, 16'hBD13, 16'hD5D7, 16'hDE59, 16'hE6DB, 16'hF75D, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'hDDD7, 16'h934D, 16'h9B4D, 16'hCD96, 16'hE659, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFF9F, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hFF1D, 16'hF69C, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEDD9, 16'hEDD9, 16'hE5D9, 16'hEDD9, 16'hDD57, 16'h9B4E, 16'hB411, 16'hEDD8, 16'hEE1A, 16'hE619, 16'hE619, 16'hE61A, 16'hE61A, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE19, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hEE5A, 16'hDD56, 16'hABCF, 16'hE5D8, 16'hEE5A, 16'hEE5A, 16'hD597, 16'hD515, 16'hDD96, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hDDD7, 16'hE5D7, 16'hE5D7, 16'hDDD7, 16'hE618,
        16'hAC10, 16'hD596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'h9A8B, 16'hCC53, 16'hF598, 16'hF5D9, 16'hDCD4, 16'hA2CB, 16'hAB4E, 16'hE597, 16'hEE1A, 16'hE5D9, 16'hE5D9, 16'hE619, 16'hE619, 16'hE619, 16'hE5D9, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619,
        16'hE61A, 16'hE619, 16'hEE19, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE19, 16'hEE1A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE61A, 16'hE5D9, 16'hE5D8, 16'hDD57, 16'hD516, 16'hD515, 16'hC493, 16'hA34D, 16'h928B, 16'hB3D0, 16'h9ACC, 16'h928A, 16'hA38D, 16'hB451, 16'hC555, 16'hEEDB, 16'hEEDB, 16'hCD96, 16'h9B4D, 16'hBC52, 16'hE65A, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFF1D, 16'hFEDC, 16'hF69C, 16'hFE9C, 16'hFEDC, 16'hFEDC, 16'hFF1D, 16'hFF5E, 16'hFF1D, 16'hF69C, 16'hFE9B, 16'hF65B, 16'hF69B, 16'hF69B, 16'hFE9B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEDD9, 16'hEDD9, 16'hE5D9, 16'hE5D8, 16'hE598, 16'hC4D4, 16'hCD15, 16'hEE19, 16'hEE1A, 16'hE619, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619,
        16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE1A, 16'hE619, 16'hB410, 16'hD556, 16'hEE19, 16'hD556, 16'hF6DC, 16'hFFDF, 16'hF71D, 16'hE65A, 16'hD596, 16'hDD96, 16'hE597, 16'hE5D8, 16'hE5D7, 16'hE5D7, 16'hE5D8, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D8, 16'hE5D7, 16'hE5D7, 16'hDDD7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D8, 16'h9B4D, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hBC11, 16'hB30D, 16'hED97, 16'hF619, 16'hFE19, 16'hED97, 16'hC3D0, 16'hAACC, 16'hD515, 16'hEE19, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE61A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE61A, 16'hE5D9, 16'hE598, 16'hE598, 16'hDD57, 16'hD556, 16'hDD56, 16'hC493, 16'h8A8A, 16'h928A,
        16'h9B0C, 16'hC514, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF1D, 16'hF6DC, 16'hF69B, 16'hFE9B, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hF69C, 16'hF69C, 16'hFE9B, 16'hF65B, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hDD57, 16'hEDD8, 16'hE5D9, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hE619, 16'hEDD9, 16'hEDD9, 16'hE5D9, 16'hEDD9, 16'hDD97, 16'hD556, 16'hE619, 16'hEE1A, 16'hE61A, 16'hE619, 16'hE61A, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE5A, 16'hEE19, 16'hCD15, 16'hDD97, 16'hEE1A, 16'hEE19, 16'hEE5A, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hEEDC, 16'hE618, 16'hDD96, 16'hE5D7, 16'hE5D7, 16'hE5D8, 16'hE5D7, 16'hE5D7, 16'hE5D7,
        16'hE5D7, 16'hE5D7, 16'hE5D8, 16'hE5D7, 16'hE5D7, 16'hDDD7, 16'hDDD7, 16'hE5D7, 16'hE5D7, 16'hDDD7, 16'hE5D8, 16'hDD97, 16'h9B0C, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDD96, 16'hBB0E, 16'hF5D8, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hFDD9, 16'hD492, 16'h99C8, 16'hBC11, 16'hEE19, 16'hEE1A, 16'hE619, 16'hE619, 16'hE619, 16'hE61A,
        16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hE619, 16'hE619, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hEE1A, 16'hE61A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE61A, 16'hEE1A, 16'hE619, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hEE1A, 16'hE5D8, 16'hBC51, 16'hC493, 16'hD5D8, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hFEDD, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9B, 16'hF69B, 16'hF65B, 16'hF65B, 16'hF61A, 16'hE598, 16'hF65A, 16'hFE9B, 16'hF65A, 16'hEE1A, 16'hEE1A, 16'hE598, 16'hE598, 16'hE5D8, 16'hE598, 16'hD516, 16'hE5D8, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hEE19, 16'hE619, 16'hE619, 16'hE619, 16'hEE1A, 16'hE61A,
        16'hE61A, 16'hE61A, 16'hEE1A, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE19, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE61A, 16'hE5D8, 16'hD555, 16'hD555, 16'hD556, 16'hE5D8, 16'hDD97, 16'hD556, 16'hEE9B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9A, 16'hE597, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hDDD7, 16'hE5D7, 16'hDDD7, 16'hE618, 16'hCD55, 16'hA34D, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9A, 16'hC30D, 16'hF597, 16'hF619, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hFDD9, 16'hE515, 16'hAB0D, 16'hBC10, 16'hE598, 16'hEE1A, 16'hE619, 16'hE619, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hEE1A, 16'hE61A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE61A, 16'hEE1A, 16'hE619, 16'hE5D9, 16'hDDD9,
        16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hEE1A, 16'hE5D8, 16'hBC52, 16'hA38E, 16'hCD56, 16'hFF5E, 16'hFFDF, 16'hFF9F, 16'hFF1D, 16'hF69B, 16'hF65A, 16'hEE19, 16'hEE19, 16'hF65B, 16'hFE9B, 16'hF65B, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE5D8, 16'hBC52, 16'hCC94, 16'hE597, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hDD57, 16'hCCD5, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hDD97, 16'hEDD9, 16'hEE19, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE619, 16'hE619, 16'hE61A, 16'hEE1A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE19, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE5D8, 16'hBC92, 16'hB411, 16'hCD14, 16'hCCD4, 16'hCCD4, 16'hEE19, 16'hF6DB, 16'hF71C, 16'hF75D,
        16'hFF5E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hDDD7, 16'hDDD7, 16'hDDD7, 16'hE618, 16'hC4D3, 16'hA38E, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hCC11, 16'hE4D4, 16'hFE19,
        16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hFE19, 16'hF598, 16'hBBCF, 16'hA2CB, 16'hDD56, 16'hEE1A, 16'hE61A, 16'hE619, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hE619, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hDDD9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE619, 16'hE5D8, 16'hCCD4, 16'h930C, 16'hBC93, 16'hF6DC, 16'hFF9F, 16'hFF5D, 16'hF69B, 16'hEE19, 16'hEE19, 16'hDD97, 16'hD515, 16'hD556, 16'hEDD9, 16'hEE1A, 16'hEE19, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hB3D0, 16'hAB8F, 16'hE5D8, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hE619, 16'hE5D9, 16'hE5D9, 16'hEDD9, 16'hCCD4, 16'hDD98, 16'hDDD8, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hD515,
        16'hC493, 16'hDD57, 16'hEDD9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE19, 16'hEE19, 16'hEE19, 16'hE619, 16'hEE1A, 16'hEE19, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE5D9, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE19, 16'hE619, 16'hEE19, 16'hEE1A, 16'hE5D8, 16'hC492, 16'hC493, 16'hD515, 16'hEE5A, 16'hFF5D, 16'hF71C, 16'hEEDB, 16'hE69A, 16'hEEDB, 16'hE69A, 16'hEEDC, 16'hF71D, 16'hF75E, 16'hFF9F, 16'hEE9B, 16'hE597, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hDDD7, 16'hE618, 16'hB451, 16'hB451, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD514, 16'hDC12, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hDCD4, 16'hAB0C, 16'hC452, 16'hEE19, 16'hEE1A, 16'hE619, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A,
        16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hDDD8, 16'hE5D8, 16'hE5D8, 16'hDDD8, 16'hE5D9, 16'hE619, 16'hCD15, 16'h8ACB, 16'h9B4E, 16'hDD97, 16'hFE9C, 16'hF69B, 16'hEE5A, 16'hE5D8, 16'hE5D8, 16'hE557, 16'hC493, 16'hC494, 16'hDD56, 16'hEE19, 16'hE619, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D9, 16'hC452, 16'hA30D, 16'hE557, 16'hEE1A, 16'hE5D9, 16'hEE19, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hDD56, 16'hDD97, 16'hE5D8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hE5D9, 16'hDD56, 16'hC452, 16'hD516, 16'hE5D8, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hD557, 16'hE5D8, 16'hEE19, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D9, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE1A, 16'hEE1A, 16'hEE1A,
        16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE19, 16'hEE19, 16'hDD97, 16'hCD15, 16'hD556, 16'hE619, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hF71C, 16'hEE9A, 16'hE659, 16'hE618, 16'hD596, 16'hCD55, 16'hDDD7, 16'hE5D7, 16'hE5D7, 16'hE5D8, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hDDD7, 16'hE618, 16'hA38E, 16'hC4D3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF69B, 16'hD390, 16'hF5D8, 16'hFE1A, 16'hF5D9, 16'hF619, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hFE19, 16'hE516, 16'hAB0C, 16'hC411, 16'hE5D8, 16'hEE1A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE619, 16'hE5D9, 16'hDDD8, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hE619, 16'hDD97, 16'hABD0, 16'h824A, 16'hC493, 16'hEE19, 16'hF65A, 16'hEDD9, 16'hE5D8, 16'hE5D8, 16'hE597, 16'hCCD4, 16'hBC53, 16'hD556, 16'hE5D8, 16'hE5D9, 16'hE5D8, 16'hDD98, 16'hDDD8, 16'hE5D8, 16'hDDD8, 16'hE5D9, 16'hCC93, 16'hA30D, 16'hD4D4, 16'hEE19, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9,
        16'hE5D9, 16'hE5D9, 16'hDD57, 16'hD556, 16'hE5D8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hE5D8, 16'hE5D8, 16'hCCD4, 16'hCCD4, 16'hDD98, 16'hE5D9, 16'hE5D8, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDDD8, 16'hDDD8, 16'hD556, 16'hC493, 16'hCD15, 16'hDD98, 16'hE5D9, 16'hE5D8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDDD8, 16'hE5D9, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE19, 16'hDD97, 16'hD556, 16'hDDD8, 16'hEE19, 16'hEE1A, 16'hEE5A, 16'hEE1A, 16'hE619, 16'hE5D9, 16'hDD57, 16'hE597, 16'hE597, 16'hDD97, 16'hD597, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hF71C, 16'hE659, 16'hE5D7, 16'hE597, 16'hE5D8, 16'hE5D8, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hA38E, 16'hD5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD492, 16'hDCD4, 16'hFE1A, 16'hF619, 16'hF619, 16'hF619, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF619, 16'hED97, 16'hC3CF, 16'hAB4D, 16'hDD15, 16'hEE1A, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE61A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE1A,
        16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE619, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hE5D9, 16'hCCD5, 16'h8A8A, 16'hA38F, 16'hDD98, 16'hEE19, 16'hE5D9, 16'hE5D8, 16'hE598, 16'hE5D8, 16'hDD56, 16'hBC52, 16'hC4D4, 16'hDD98, 16'hE5D9, 16'hE5D8, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hE5D8, 16'hD516, 16'hB38E, 16'hBBD0, 16'hED98, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hE598, 16'hD556, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hE5D9, 16'hDD97, 16'hB411, 16'hCD15, 16'hE5D9, 16'hE5D8, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hDDD8, 16'hE5D8, 16'hDD97, 16'hCCD4, 16'hBC52, 16'hD516, 16'hE5D8, 16'hDDD8, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hE5D9, 16'hE619, 16'hE619,
        16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hCD15, 16'hB452, 16'hABD0, 16'hB451, 16'hC493, 16'hCD15, 16'hE5D8, 16'hEE5A, 16'hD597, 16'hCD15, 16'hD515, 16'hC493, 16'hDDD8, 16'hE618, 16'hDD97, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5D, 16'hEE59, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D8, 16'hDDD7, 16'hAB8E, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE597, 16'hD3D0, 16'hF619, 16'hF619, 16'hF619, 16'hF619, 16'hF619, 16'hF619, 16'hF619, 16'hF619, 16'hF5D9, 16'hFE19, 16'hF5D8, 16'hD492, 16'h9249, 16'hCCD3, 16'hEE5A, 16'hEE1A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hE61A, 16'hE61A, 16'hE619, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hE5D9, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hE5D8, 16'hDD97, 16'hA38F, 16'h8A8B, 16'hC493, 16'hEDD9, 16'hE5D9, 16'hE5D8, 16'hDD98, 16'hDD98, 16'hE5D8, 16'hCD15, 16'hB411, 16'hD516, 16'hE5D9, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hDD98,
        16'hDD98, 16'hBC11, 16'hB38F, 16'hD4D4, 16'hE5D9, 16'hE5D8, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hE5D9, 16'hE5D8, 16'hDD57, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hE5D9, 16'hDD98, 16'hBC52, 16'hCCD4, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hE5D8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hE5D8, 16'hDD57, 16'hCCD4, 16'hD515, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hE5D9, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE19, 16'hEE19, 16'hE5D8, 16'hDD97, 16'hD556, 16'hBC51, 16'h930C, 16'hDD97, 16'hEE1A, 16'hE619, 16'hEE19, 16'hEE5A, 16'hE65A, 16'hE65A, 16'hE618, 16'hD556, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hEEDB, 16'hDE18, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hDDD7, 16'hDDD7, 16'hDDD7, 16'hDDD7,
        16'hDDD7, 16'hDE18, 16'hCD55, 16'hA3CF, 16'hFF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF69B, 16'hD38F, 16'hF5D8, 16'hFE1A, 16'hF619, 16'hF619, 16'hF619, 16'hF619, 16'hF619, 16'hF619, 16'hF619, 16'hF5D9, 16'hF5D9, 16'hF5D8, 16'hDD15, 16'hAB4D, 16'hA38E, 16'hE5D9, 16'hEE5A, 16'hE61A, 16'hEE1A, 16'hE61A,
        16'hE619, 16'hEE19, 16'hEE1A, 16'hE61A, 16'hE61A, 16'hE619, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE5D9, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDDD8, 16'hDD97, 16'h9B0D, 16'hA34E, 16'hDD97, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hDDD8, 16'hDD98, 16'hE598, 16'hC493, 16'hBC52, 16'hDD97, 16'hE5D8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD97, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hE5D8, 16'hD516, 16'hC411, 16'hC452, 16'hDD97, 16'hE5D8, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDD97, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDD98, 16'hC494, 16'hCD15, 16'hE5D8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hE5D8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDD98,
        16'hDD98, 16'hDD98, 16'hE5D8, 16'hDD56, 16'hCCD5, 16'hD556, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDDD8, 16'hE5D9, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE1A, 16'hEE1A, 16'hDD97, 16'hC493, 16'hC4D3, 16'hCD15, 16'hE619, 16'hEE5A, 16'hDDD8, 16'hCD15, 16'hDDD8, 16'hE619, 16'hDDD8, 16'hE619, 16'hD556, 16'hE659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'hDDD7, 16'hDDD7, 16'hE5D7, 16'hE5D7, 16'hE5D7, 16'hDDD7, 16'hDDD7, 16'hDDD7, 16'hDDD8, 16'hDE19, 16'hB492, 16'hB451, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hDC93, 16'hE514, 16'hFE5A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF619, 16'hF619, 16'hF619, 16'hF619, 16'hF619, 16'hF5D9, 16'hF5D9, 16'hF619, 16'hE556, 16'hAB4E, 16'hA30D, 16'hDD97, 16'hEE5A, 16'hE61A, 16'hEE1A, 16'hE61A, 16'hE61A, 16'hEE19, 16'hE619, 16'hE61A, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hE619, 16'hE5D9, 16'hDDD8, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hE5D8, 16'hD556, 16'h92CB, 16'hBC52, 16'hEDD9, 16'hE5D9, 16'hE598, 16'hDD98, 16'hDD98, 16'hE598, 16'hE598, 16'hC452, 16'hC493,
        16'hE5D8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hC494, 16'hC493, 16'hCCD5, 16'hE5D8, 16'hDD98, 16'hE5D8, 16'hDDD8, 16'hDDD8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE5D8, 16'hE598, 16'hDD97, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDD98, 16'hDDD8, 16'hE5D9, 16'hC494, 16'hCCD4, 16'hE5D8, 16'hDD98, 16'hDDD8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDDD8, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hE5D8, 16'hDD97, 16'hCCD5, 16'hCCD5, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hEE1A, 16'hEE19, 16'hD556, 16'hC492, 16'hB411, 16'hCD15, 16'hEE5A, 16'hEE9B, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hCD56, 16'hDDD7, 16'hFF5E, 16'hF75D, 16'hF75E, 16'hFF9E, 16'hF79D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE659, 16'hDD97, 16'hDDD7, 16'hDDD7, 16'hDDD7, 16'hDDD7, 16'hDDD7, 16'hDDD8, 16'hDDD8, 16'hDE19, 16'hAC10, 16'hCD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE18, 16'hD3D0, 16'hF619, 16'hFE1A, 16'hFE1A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF619,
        16'hF619, 16'hF619, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF619, 16'hF5D8, 16'hBC10, 16'h924A, 16'hDD56, 16'hEE5A, 16'hEE1A, 16'hE61A, 16'hE61A, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE5D9, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hE5D8, 16'hCCD4, 16'h8ACC, 16'hD515, 16'hEE1A, 16'hE5D8, 16'hE598, 16'hE598, 16'hE598, 16'hE5D8, 16'hDD57, 16'hB3D0, 16'hC493, 16'hE5D9, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD97, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD57, 16'hBC52, 16'hC493, 16'hDD97, 16'hDD98, 16'hE598, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hDD98, 16'hDD57, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hE5D8,
        16'hC493, 16'hD516, 16'hE5D9, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hE598, 16'hCD15, 16'hC4D4, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hE5D9, 16'hE619, 16'hE619, 16'hE619, 16'hEE1A, 16'hE619, 16'hD556, 16'hABD0, 16'h9B8E, 16'hD557, 16'hF69B, 16'hF69B, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hDD97, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hE5D8, 16'hDDD7, 16'hDDD7, 16'hDDD7, 16'hDDD7, 16'hDDD8, 16'hDDD8, 16'hDE18, 16'hD5D8, 16'h9B4D, 16'hE658, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFEDC, 16'hF69C, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'hCBD0, 16'hED57, 16'hFE5B, 16'hF65A, 16'hFE1A, 16'hFE1A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF619, 16'hF619, 16'hF619, 16'hF619, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hC451, 16'h9249, 16'hDD56, 16'hEE1A, 16'hE61A, 16'hEE19, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE61A, 16'hEE19, 16'hE619, 16'hE5D8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hE5D8, 16'hC4D4, 16'hA34E,
        16'hE598, 16'hF65A, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDD97, 16'hB3D0, 16'hCCD4, 16'hE5D9, 16'hDD98, 16'hDDD8, 16'hE5D8, 16'hDDD8, 16'hDD98, 16'hDD97, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hD556, 16'hC493, 16'hD515, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hDD97, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hE598, 16'hC493, 16'hD516, 16'hE5D9, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hE5D8, 16'hCCD5, 16'hC494, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hE5D9, 16'hEE19, 16'hE619, 16'hCD15, 16'hAC10, 16'hC4D3, 16'hCD15, 16'hE5D9, 16'hE619, 16'hDD97, 16'hE619, 16'hF65B, 16'hEE9B, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5B,
        16'hEE5B, 16'hCD56, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hF75E, 16'hFF5E, 16'hE69A, 16'hEEDB, 16'hF75D, 16'hFF9E, 16'hFFDF, 16'hFF9E, 16'hF75D, 16'hEE9B, 16'hDDD7, 16'hDDD7, 16'hDDD7, 16'hDDD8, 16'hDE18, 16'hDE18, 16'hDE19, 16'hCD56, 16'hA38E, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF1D, 16'hF6DC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDCD4, 16'hE4D4, 16'hFE5B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF619, 16'hF619, 16'hF619, 16'hF5D9, 16'hF619, 16'hF619, 16'hCC93, 16'h9289, 16'hCCD4, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE5D9, 16'hE5D8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDD98, 16'hE5D9, 16'hCCD4, 16'hAB8E, 16'hEDD9, 16'hFE9B, 16'hEE1A, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hE598, 16'hB411, 16'hCCD5, 16'hE5D9, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD97, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hE5D8, 16'hD515, 16'hCC93, 16'hD557, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE5D8, 16'hDD98, 16'hDD98, 16'hE5D8, 16'hDDD8,
        16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDDD8, 16'hDD97, 16'hC453, 16'hDD97, 16'hE598, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hCCD5, 16'hC493, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hE5D8, 16'hD556, 16'hB452, 16'hBC93, 16'hD556, 16'hEE5A, 16'hEE1A, 16'hE61A, 16'hDD98, 16'hBC52, 16'hBC92, 16'hCD14, 16'hD597, 16'hE619, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hCD15, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hEEDB, 16'hEEDB, 16'hEE9A, 16'hD618, 16'hD5D7, 16'hDE18, 16'hEEDB, 16'hF6DC, 16'hCD55, 16'hE619, 16'hDE19, 16'hD5D8, 16'hDE18, 16'hDE18, 16'hDE18, 16'hD618, 16'hDE59, 16'hBCD3, 16'hABCF, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE59, 16'hD3D0, 16'hF61A, 16'hFE5B, 16'hFE5A, 16'hFE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF619, 16'hF619, 16'hF619, 16'hF619, 16'hFE1A, 16'hDD15, 16'h9ACB, 16'hCC94, 16'hEE1A, 16'hE61A, 16'hE619, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hE5D9, 16'hE5D8,
        16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hE5D8, 16'hCD15, 16'hBC10, 16'hF65A, 16'hF69B, 16'hF65B, 16'hF69B, 16'hEE1A, 16'hE5D9, 16'hE5D9, 16'hE598, 16'hC452, 16'hCCD4, 16'hE5D9, 16'hDD98, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDDD8, 16'hDD97, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDD98, 16'hE5D8, 16'hCCD5, 16'hCCD4, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hDD97, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE5D8, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hE5D9, 16'hD556, 16'hC494, 16'hE598, 16'hDD98, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hE5D8, 16'hC494, 16'hBC53, 16'hE598, 16'hDD98, 16'hDD98, 16'hDD98, 16'hE5D8, 16'hD557, 16'hDD97, 16'hE61A, 16'hE61A,
        16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE5D8, 16'hDD56, 16'hBC51, 16'h92CB, 16'hA38E, 16'hE5D8, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE9B, 16'hE619, 16'hCD56, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'hEEDB, 16'hEEDB, 16'hEEDB, 16'hEEDC, 16'hEEDB, 16'hDE18, 16'hCD55, 16'hD5D7, 16'hE659, 16'hE65A, 16'hD5D8, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hDE19, 16'hA3CF, 16'hCD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5D, 16'hD451, 16'hED56, 16'hFE9B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF619, 16'hF619, 16'hF619, 16'hF619, 16'hF61A, 16'hDD56, 16'h928A, 16'hC493, 16'hEE1A, 16'hE61A, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE5D9, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hE5D8, 16'hDD57, 16'hC412, 16'hEE19, 16'hF65A, 16'hEE19, 16'hF69C, 16'hFEDD, 16'hF65B, 16'hEDD9, 16'hE5D9, 16'hD4D4, 16'hCCD4, 16'hE5D9, 16'hDD98, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDD98, 16'hDD97, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDD98, 16'hE5D8, 16'hD516, 16'hCCD5, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hE5D8, 16'hE5D8, 16'hE5D8,
        16'hE5D8, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hDD98, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hE5D9, 16'hCCD4, 16'hD515, 16'hE598, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hB3D1, 16'hCCD4, 16'hDDD8, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hE619, 16'hE619, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE619, 16'hE619, 16'hCD56, 16'hAC11, 16'hB451, 16'hCCD4, 16'hDD97, 16'hD515, 16'hDD97, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE9B, 16'hDDD8, 16'hE69A, 16'hFFDF, 16'hFF9E, 16'hF71C, 16'hEEDB, 16'hEEDB, 16'hEE9B, 16'hEEDB, 16'hEEDB, 16'hF71C, 16'hF6DB, 16'hE659, 16'hCD97, 16'hD5D8, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD5D7, 16'h9B4D, 16'hEE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDD95, 16'hD452, 16'hFE5B, 16'hF65B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hFE5A, 16'hFE5A, 16'hF65A, 16'hF61A, 16'hF61A, 16'hF619, 16'hF619, 16'hF65A, 16'hE597, 16'hA2CC, 16'hBC12, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hEE1A, 16'hEE1A,
        16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE619, 16'hEE19, 16'hE619, 16'hE5D8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDDD8, 16'hDD57, 16'hCC53, 16'hED99, 16'hEDD8, 16'hCC11, 16'hF65B, 16'hFF5E, 16'hF6DC, 16'hEE1A, 16'hEDD9, 16'hE556, 16'hCC93, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hE5D8, 16'hDD97, 16'hD557, 16'hE598, 16'hDD98, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hDD98, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hCCD4, 16'hD556, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98,
        16'hDD98, 16'hDD98, 16'hDD97, 16'hB411, 16'hD556, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDDD9, 16'hDDD9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hDDD8, 16'hE5D9, 16'hEDD9, 16'hDD97, 16'hBC92, 16'hB451, 16'hE619, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hDE19, 16'hF71D, 16'hFFDF, 16'hF71C, 16'hEEDB, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEEDB, 16'hEEDC, 16'hF71C, 16'hEEDB, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hDE19, 16'hC555, 16'hAC0F, 16'hFF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF6DB, 16'hCB8F, 16'hF5D8, 16'hFE9B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hF65A, 16'hF65A, 16'hF61A, 16'hFE5A, 16'hF61A, 16'hEDD9, 16'hF61A, 16'hE5D8, 16'hA2CC, 16'hB411, 16'hEE19, 16'hEE1A, 16'hE619, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hE5D8, 16'hCC53, 16'hE557, 16'hED57, 16'hD411, 16'hF69B, 16'hFF5E, 16'hF6DD, 16'hF65B, 16'hF61A, 16'hF5D9, 16'hD4D4, 16'hED98, 16'hE599, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hDD98, 16'hE598, 16'hDD98, 16'hDDD8, 16'hE5D8, 16'hDDD8,
        16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE598, 16'hE5D8, 16'hDD98, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDDD8, 16'hDD97, 16'hD515, 16'hDD57, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hE5D8, 16'hCD15, 16'hBC52, 16'hDD98, 16'hDD97, 16'hDD98, 16'hDDD8, 16'hDDD9, 16'hDDD9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE619, 16'hD556, 16'hB451, 16'hB452, 16'hD556, 16'hEE5A, 16'hEE9B, 16'hE65A, 16'hE65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hE619, 16'hDE59, 16'hFF9E, 16'hFF9E, 16'hEEDB, 16'hEE9B, 16'hE69A, 16'hEE9B, 16'hEE9B, 16'hE69A, 16'hEEDB, 16'hF6DC, 16'hF6DC, 16'hEE9B, 16'hD618, 16'hD618,
        16'hD618, 16'hD618, 16'hD618, 16'hDE19, 16'hA451, 16'hBC92, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hD4D3, 16'hE4D5, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE9B, 16'hFE9B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hF65B,
        16'hF61A, 16'hDD57, 16'hCC94, 16'hD515, 16'hE5D8, 16'hF69B, 16'hEDD8, 16'hA30D, 16'hB3D0, 16'hE5D8, 16'hEE1A, 16'hE619, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hEE19, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hE5D8, 16'hCC93, 16'hE557, 16'hED57, 16'hD452, 16'hFEDC, 16'hFF9F, 16'hF6DD, 16'hF65B, 16'hF65B, 16'hF61A, 16'hDD15, 16'hE597, 16'hEDD9, 16'hE5D8, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDD98, 16'hDD98, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hDD57, 16'hDD98, 16'hDD98, 16'hDD98, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hDD98, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDDD8, 16'hDD98, 16'hE598, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hE598, 16'hD515, 16'hD516, 16'hD557,
        16'hDD97, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hE5D8, 16'hBC52, 16'hC4D4, 16'hDD97, 16'hDD97, 16'hDDD8, 16'hDDD9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hD556, 16'hCD16, 16'hE5D8, 16'hE5D8, 16'hD596, 16'hE619, 16'hEE5A, 16'hE65A, 16'hE619, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE619, 16'hE69A, 16'hF75D, 16'hEEDC, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE69A, 16'hD618, 16'hDE59, 16'hEEDB, 16'hE69A, 16'hD618, 16'hD5D8, 16'hD5D8, 16'hD618, 16'hD618, 16'hD618, 16'h8B4C, 16'hDE17, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE19, 16'hD3D1, 16'hF65A, 16'hFE9B, 16'hFE5B, 16'hFE9B, 16'hFE9B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hCCD4, 16'hCC92, 16'hEDD8, 16'hF69B, 16'hF69B, 16'hEE5A, 16'hF65A, 16'hEE19, 16'hB3D0, 16'hA38F, 16'hE5D8, 16'hEE1A, 16'hE619, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hE619, 16'hE619, 16'hE5D9, 16'hE5D9, 16'hDDD8, 16'hDD98, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hE5D8, 16'hD4D4, 16'hDCD5, 16'hED98, 16'hCC52, 16'hFF1D, 16'hFFDF, 16'hFF5E, 16'hF65B, 16'hF65B, 16'hFE5B, 16'hE556, 16'hE556, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hE5D9,
        16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDD98, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hCCD4, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hDD98, 16'hE5D8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD97, 16'hD4D5, 16'hD516, 16'hCCD4, 16'hDD98, 16'hDD97, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hD557, 16'hB412, 16'hD556, 16'hDD57, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hE5D8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hD597, 16'hCD15, 16'hBC52, 16'hB451, 16'hBC93, 16'hDDD8, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE65A, 16'hE65A, 16'hDE19, 16'hEEDB,
        16'hEEDB, 16'hEE9A, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE69A, 16'hDE18, 16'hD5D7, 16'hD618, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD618, 16'hDE59, 16'hBD14, 16'h8B0C, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF1D, 16'hD411,
        16'hED98, 16'hFE9C, 16'hF65B, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE5B, 16'hFE5B, 16'hFE9B, 16'hEDD8, 16'hDD56, 16'hDD56, 16'hCD15, 16'hD515, 16'hEE1A, 16'hEE5A, 16'hF69B, 16'hF65A, 16'hB390, 16'h9B0C, 16'hDD57, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hE619, 16'hE5D9, 16'hE5D8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hE5D8, 16'hDD16, 16'hDCD5, 16'hED58, 16'hCC11, 16'hFF1D, 16'hFFDF, 16'hFF9E, 16'hF6DC, 16'hF65B, 16'hFE5B, 16'hED98, 16'hDCD4, 16'hF61A, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE598, 16'hE5D8, 16'hDD97, 16'hD4D4, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hDD97, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8,
        16'hE5D8, 16'hDD98, 16'hE5D8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hE5D8, 16'hD516, 16'hD516, 16'hCCD5, 16'hCCD5, 16'hDD57, 16'hD556, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD97, 16'hDD98, 16'hC4D4, 16'hBC52, 16'hDD57, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hD597, 16'hDD97, 16'hD597, 16'hD597, 16'hD557, 16'hD557, 16'hD557, 16'hD597, 16'hDD97, 16'hD597, 16'hBC93, 16'hAC11, 16'hC4D4, 16'hDDD8, 16'hDDD9, 16'hDE19, 16'hE659, 16'hE65A, 16'hDE18, 16'hE65A, 16'hEE9B, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE69A, 16'hDE19, 16'hD5D7, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD618, 16'hDE19, 16'h9C10, 16'hB4D3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDD15, 16'hDC94, 16'hFE9C, 16'hF69B, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE5B, 16'hFE9B, 16'hFE9B, 16'hF65A, 16'hEE19, 16'hE5D8, 16'hEE19, 16'hEE19, 16'hDDD8, 16'hE5D8, 16'hF69A, 16'hC4D3, 16'hA30C, 16'hCCD4, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDDD8, 16'hE5D8, 16'hE597, 16'hD494, 16'hED98, 16'hCC12, 16'hF69B, 16'hFFDF,
        16'hFF9F, 16'hF6DD, 16'hF69B, 16'hFE9C, 16'hF61A, 16'hDC95, 16'hF5D9, 16'hF61A, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hE5D9, 16'hE598, 16'hE5D8, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE5D9, 16'hDD16, 16'hDD16, 16'hE5D9, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDD97, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hC494, 16'hDD57, 16'hC4D4, 16'hD516, 16'hD516, 16'hD516, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hD556, 16'hA390, 16'hC4D4, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD16, 16'hD556, 16'hD556, 16'hD557, 16'hD557,
        16'hD557, 16'hD597, 16'hDD98, 16'hD556, 16'hBC93, 16'hBC93, 16'hD597, 16'hDDD8, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE65A, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE65A, 16'hE69A, 16'hE65A, 16'hDE19, 16'hD5D7, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD619, 16'hCDD7, 16'h8B4D, 16'hDE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF65A, 16'hCBD0, 16'hF61A, 16'hFE9C, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hF69B, 16'hF65A, 16'hEE19, 16'hE5D8, 16'hE619, 16'hDDD7, 16'hE619, 16'hEEDC, 16'hF75E, 16'hFFDF, 16'hFF5E, 16'hDD97, 16'hB411, 16'hE5D8, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hC452, 16'hDD16, 16'hD453, 16'hE5D9, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hF69C, 16'hF69C, 16'hFE5B, 16'hE495, 16'hEDD9, 16'hFE5B, 16'hF61A, 16'hF61A, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hE598, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE5D9, 16'hD4D4, 16'hDD57, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8,
        16'hE5D8, 16'hE5D8, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hE5D8, 16'hD516, 16'hCCD4, 16'hDD97, 16'hC493, 16'hDD57, 16'hCCD5, 16'hDD57, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD97, 16'hD597, 16'hDD57, 16'hC4D4, 16'hA38F, 16'hCD15, 16'hD516, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD16, 16'hC515, 16'hD556, 16'hCD56, 16'hD556, 16'hD556, 16'hD557, 16'hCD16, 16'hCD15, 16'hCD14, 16'hC4D4, 16'hBC92, 16'hC4D4, 16'hD597, 16'hD5D8, 16'hD5D8, 16'hDE19, 16'hDE59, 16'hE659, 16'hE65A, 16'hDE59, 16'hDE59, 16'hDE59, 16'hDE19, 16'hD5D8, 16'hCDD7, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD618, 16'hD618, 16'hD619, 16'hACD3, 16'h9C10, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD493, 16'hE516, 16'hFE9C, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE9C, 16'hF65A, 16'hDD56, 16'hE618, 16'hE659, 16'hEEDB, 16'hF75D, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hF6DC, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE5A, 16'hEE1A, 16'hE5D9, 16'hE5D9,
        16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D9, 16'hDD16, 16'hDCD5, 16'hDC94, 16'hDD56, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFEDD, 16'hFEDD, 16'hFEDD, 16'hED98, 16'hED16, 16'hFE5B, 16'hF65B, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF5DA, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hE598, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D9, 16'hED98, 16'hCC94, 16'hE597, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDD98, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hE598, 16'hCCD4, 16'hDD57, 16'hD516, 16'hC494, 16'hDD57, 16'hCCD4, 16'hDD97, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hD557, 16'hD556, 16'hCD16, 16'hD516, 16'hA390,
        16'hBC52, 16'hC4D4, 16'hCD16, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hD556, 16'hC4D4, 16'hA38F, 16'hABD0, 16'hABCF, 16'hBC92, 16'hB452, 16'hD597, 16'hD5D8, 16'hD597, 16'hCD56, 16'hDDD8, 16'hDE19, 16'hDE59, 16'hDE59, 16'hDE19, 16'hD5D8, 16'hD5D7, 16'hCDD7, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD619, 16'hBD55, 16'h6A8A, 16'h72CA, 16'h9C51, 16'hC5D7, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE19, 16'hD452, 16'hFE5B, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9B, 16'hFE9C, 16'hFEDC, 16'hF65A, 16'hCCD3, 16'hDD56, 16'hEE5A, 16'hF6DC, 16'hEEDC, 16'hEEDB, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hF69B, 16'hEE19, 16'hEE1A, 16'hF71D, 16'hFF9F, 16'hFF5D, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hD494, 16'hE516, 16'hD4D4, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF1E, 16'hFF1D, 16'hFF1E, 16'hF65B, 16'hE4D5, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF5D9, 16'hF61A, 16'hE598, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hEDD9, 16'hE598, 16'hCC93, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8,
        16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hE5D8, 16'hDD56, 16'hCCD4, 16'hE598, 16'hCCD4, 16'hD515, 16'hD515, 16'hCCD4, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hD597, 16'hD556, 16'hCD16, 16'hCD16, 16'hCD16, 16'hBC93, 16'hABD0, 16'hC493, 16'hC4D5, 16'hCD56, 16'hCD16, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hD557, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hBCD3, 16'hAC51, 16'hA3D0, 16'h9B8F, 16'hCD15, 16'hD597, 16'hD597, 16'hCD56, 16'hC515, 16'hDE18, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D7, 16'hCD97, 16'hCDD7, 16'hCDD8, 16'hCDD8, 16'hD5D8, 16'hD5D8, 16'hCDD8, 16'hD618, 16'hCDD8, 16'hCDD8, 16'hCDD7, 16'hAC91, 16'h58C0, 16'h9410, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'hD411, 16'hF619, 16'hFEDC, 16'hFE9C, 16'hFE9C, 16'hFE9B, 16'hFEDC, 16'hF69B, 16'hDD96, 16'hD514, 16'hEE19, 16'hE5D8, 16'hE5D8, 16'hDDD7, 16'hDD97, 16'hDDD8, 16'hEEDB, 16'hFFDF, 16'hFFDF,
        16'hFF9E, 16'hF75D, 16'hE65A, 16'hDD97, 16'hD515, 16'hE5D9, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hF6DC, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D9, 16'hD494, 16'hE516, 16'hD493, 16'hFF1D, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5F, 16'hFF1E, 16'hE516, 16'hED99, 16'hFE9C, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE1A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hE598, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hE557, 16'hCC93, 16'hE5D8, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hCCD4, 16'hDD56, 16'hDD57, 16'hC494, 16'hDD57, 16'hCCD4, 16'hD516,
        16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD97, 16'hD557, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15, 16'hABD0, 16'hBC52, 16'hB452, 16'hCD16, 16'hCD16, 16'hCD56, 16'hCD56, 16'hCD16, 16'hCD56, 16'hD556, 16'hBC94, 16'hC515, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC515, 16'hBCD4, 16'hCD56, 16'hCD56, 16'hCD97, 16'hD597, 16'hC555, 16'hCD96, 16'hD5D7, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCDD7, 16'hCDD8, 16'hCDD8, 16'hD5D8, 16'hCDD8, 16'hCDD8, 16'hD618, 16'hD659, 16'hCDD8, 16'hA492, 16'h93CE, 16'hC5D7, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD514, 16'hDD15, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFEDC, 16'hEE5A, 16'hCCD3, 16'hD515, 16'hFE9B, 16'hFEDC, 16'hFEDC, 16'hFF1D, 16'hFF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hD596, 16'hBC52, 16'hCC94, 16'hDD15, 16'hEE9B, 16'hFF5E, 16'hF75D, 16'hF69B, 16'hE619, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hEE19, 16'hDD15, 16'hDCD5, 16'hDC54, 16'hE61A, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hF61B, 16'hED16, 16'hFE9C, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hF61A, 16'hF65B, 16'hEDD9, 16'hED98, 16'hF61A, 16'hF5D9, 16'hF619, 16'hEDD9,
        16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hDD16, 16'hCC53, 16'hEDD9, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D9, 16'hE598, 16'hDD97, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hE598, 16'hDD57, 16'hD515, 16'hDD98, 16'hCCD5, 16'hCD15, 16'hDD57, 16'hC493, 16'hDD57, 16'hDD98, 16'hDD97, 16'hDD98, 16'hDD98, 16'hDD97, 16'hD556, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hCD15, 16'hBC52, 16'hABCF, 16'hB411, 16'hBC93, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD56, 16'hCD56, 16'h8B4D, 16'h7249, 16'h7A8A, 16'h9BCF, 16'hC555, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD57, 16'hCD97, 16'hCD97, 16'hC556, 16'hCD96, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97,
        16'hCDD7, 16'hCDD7, 16'hCDD8, 16'hD618, 16'hCDD8, 16'h9C51, 16'h72CB, 16'hB554, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE5A, 16'hD452, 16'hFE5B, 16'hFEDC, 16'hFEDC, 16'hF69C, 16'hD515,
        16'hE618, 16'hFEDD, 16'hFEDC, 16'hF6DC, 16'hFF1D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hF71C, 16'hF6DC, 16'hEE19, 16'hC4D4, 16'hCCD4, 16'hEDD9, 16'hE619, 16'hE5D9, 16'hE5D8, 16'hE5D9, 16'hE619, 16'hE5D8, 16'hD4D4, 16'hDD16, 16'hD556, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF1E, 16'hED57, 16'hF61B, 16'hFE9C, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hF61A, 16'hED57, 16'hF5D9, 16'hFE1A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF619, 16'hF5D9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hDD15, 16'hCC94, 16'hEDD9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hDD98, 16'hE598, 16'hDD97,
        16'hE5D8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hD515, 16'hDD57, 16'hDD57, 16'hC493, 16'hDD57, 16'hCCD5, 16'hCCD4, 16'hDD98, 16'hDD97, 16'hDD97, 16'hD597, 16'hD557, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'h9B8F, 16'hBC52, 16'hB411, 16'hCD16, 16'hCD16, 16'hCD16, 16'hD556, 16'hA3D0, 16'h71C7, 16'hBC11, 16'hC451, 16'h9B4D, 16'h8B0D, 16'hCD15, 16'hC556, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD97, 16'hCD56, 16'hCD56, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCDD7, 16'hD5D8, 16'hD618, 16'hB514, 16'h834D, 16'h9C10, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hD493, 16'hE597, 16'hFEDD, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hFEDD, 16'hFEDC, 16'hFF1D, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hF69B, 16'hF65B, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hE5D8, 16'hD556, 16'hE5D9, 16'hE619, 16'hEE1A, 16'hD4D5, 16'hE516, 16'hD4D5, 16'hFF5E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF1F, 16'hF61A, 16'hEDD8, 16'hFEDD, 16'hFE5B, 16'hF65B, 16'hF69B, 16'hFE5B, 16'hFE5B,
        16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hF619, 16'hE556, 16'hFE1B, 16'hF61A, 16'hF61A, 16'hF61A, 16'hFE1A, 16'hFE1A, 16'hF61A, 16'hF61A, 16'hF5D9, 16'hF61A, 16'hD4D5, 16'hD4D5, 16'hEDD9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDD98, 16'hE598, 16'hE598, 16'hE5D8, 16'hDD98, 16'hE5D8, 16'hEE5A, 16'hEE9B, 16'hFF1D, 16'hE5D8, 16'hE598, 16'hE598, 16'hE598, 16'hD556, 16'hD516, 16'hE598, 16'hD515, 16'hC494, 16'hDD57, 16'hC453, 16'hD516, 16'hDD97, 16'hD557, 16'hD556, 16'hD556, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hC4D5, 16'hC4D4, 16'hCD15, 16'hAC11, 16'hABCF, 16'hB411, 16'hC493, 16'hCD56, 16'hCD16, 16'hD556, 16'h828A, 16'hA38E, 16'hD493, 16'hCC92, 16'hC451, 16'h8249, 16'hAC11, 16'hD597, 16'hC514, 16'h938E, 16'hA3D0, 16'hAC51,
        16'hC515, 16'hCD97, 16'hC556, 16'hCD57, 16'hCD57, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCDD7, 16'hD5D7, 16'hBD55, 16'h9C11, 16'h93CF, 16'hA451, 16'hB4D3, 16'hBD55, 16'hAD13, 16'hEF5C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE59, 16'hD493, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hFF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hF69B, 16'hEE5A, 16'hEE5A, 16'hF65B, 16'hEE19, 16'hCD14, 16'hCCD4, 16'hE5D9, 16'hEE19, 16'hEE1A, 16'hE557, 16'hD494, 16'hDCD5, 16'hEE9B, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFEDD, 16'hE557, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFEDD, 16'hFF1D, 16'hFE9C, 16'hF65B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hED98, 16'hED98, 16'hFE5B, 16'hF61A, 16'hFE1B, 16'hFE1B, 16'hF61A, 16'hF61A, 16'hFE1A, 16'hF61A, 16'hF61A, 16'hFE1A, 16'hDCD5, 16'hE516, 16'hF619, 16'hEDD9, 16'hEDD9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDD97, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8,
        16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hEE5A, 16'hFF1D, 16'hEE19, 16'hDD98, 16'hDD98, 16'hE619, 16'hFF9F, 16'hF71D, 16'hF71D, 16'hEE5A, 16'hDD57, 16'hE598, 16'hDD97, 16'hDD97, 16'hCCD5, 16'hDD57, 16'hDD97, 16'hBC53, 16'hD516, 16'hCCD5, 16'hC453, 16'hDD57, 16'hD557, 16'hD556, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hC4D4, 16'h9B4E, 16'hB411, 16'hABD0, 16'hCD15, 16'hCD56, 16'hC4D4, 16'h7A49, 16'hC452, 16'hCC92, 16'hCC52, 16'hCC52, 16'hA30C, 16'h9B8E, 16'hCD14, 16'h7A8A, 16'h930C, 16'hA38D, 16'h8B0B, 16'h7ACB, 16'hC515, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC596, 16'hCD97, 16'hCD97, 16'hCD97, 16'hC555, 16'hAC93, 16'h9C11, 16'h834E, 16'h834D, 16'h7B4C, 16'h7B4C, 16'h6A89, 16'h9450, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hD4D4, 16'hEE19, 16'hFF1C, 16'hFEDC, 16'hFEDC, 16'hFF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5D, 16'hF69B, 16'hF65A, 16'hF69B, 16'hEE5A, 16'hD515, 16'hC492, 16'hDD56, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hEDD9, 16'hD4D4, 16'hE516, 16'hDD97, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF5F, 16'hFF5E, 16'hED98, 16'hEDD9, 16'hFEDD, 16'hF69B, 16'hF69C, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hF69C, 16'hF65B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hE556, 16'hF5D9, 16'hFE5B, 16'hFE1A, 16'hFE1B, 16'hFE1B, 16'hFE1B, 16'hF65B, 16'hFE1A, 16'hFE1A, 16'hF61A, 16'hFE5B, 16'hDC94, 16'hE516, 16'hF61A, 16'hF5D9, 16'hF5D9, 16'hEDD9, 16'hEDD9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDD57, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE65A, 16'hFF5E, 16'hFF5D, 16'hFFDF, 16'hF71D, 16'hDD98, 16'hE598, 16'hDD98, 16'hEEDC, 16'hF71D, 16'hE5D8, 16'hE5D8, 16'hDD98, 16'hDD98, 16'hDD97, 16'hE598, 16'hD516, 16'hCD15, 16'hDD98, 16'hCD15, 16'hBC52, 16'hDD56, 16'hB411, 16'hCD15, 16'hDD57, 16'hD556, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hC4D4, 16'hCCD5, 16'hA3D0, 16'hB411, 16'hB3D0, 16'hC4D4, 16'hD556, 16'hB452,
        16'h828A, 16'hCC92, 16'hCC92, 16'hCC52, 16'hCC92, 16'hB3CF, 16'h9B4D, 16'h8B0C, 16'h9B8D, 16'hABCF, 16'h6186, 16'hBC51, 16'h930C, 16'h8B4E, 16'hCD56, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hCD97, 16'hC556, 16'hC556, 16'hBD15, 16'h9C11, 16'h9C11, 16'h9410, 16'hA492, 16'h9C51, 16'h7B4C, 16'h9410, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDD97, 16'hDCD5, 16'hFEDC, 16'hFEDC, 16'hFF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFF5D, 16'hF69B, 16'hF69B, 16'hF69B, 16'hE5D8, 16'hC492, 16'hD515, 16'hEE1A, 16'hF65A, 16'hEE1A, 16'hEE19, 16'hEE5A, 16'hD515, 16'hDD57, 16'hDD16, 16'hFF1D, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hF69C, 16'hE556, 16'hFE9C, 16'hFE9B, 16'hFE5B, 16'hFE9B, 16'hFE9C, 16'hFEDD, 16'hFEDD, 16'hF65B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hF61A, 16'hE515, 16'hF61A, 16'hF65B, 16'hFE1B, 16'hFE1A, 16'hFE1A, 16'hFE5B, 16'hF61B, 16'hFE1A, 16'hFE1A, 16'hF61A, 16'hFE5B, 16'hDC94, 16'hED57, 16'hF61A, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hEDD9, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8,
        16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hCC93, 16'hDD57, 16'hE5D8, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDD98, 16'hEE9A, 16'hFFDF, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hE5D9, 16'hE598, 16'hE5D8, 16'hE598, 16'hE598, 16'hE598, 16'hDD98, 16'hE598, 16'hDD98, 16'hDD97, 16'hDD97, 16'hDD57, 16'hCCD5, 16'hDD57, 16'hDD57, 16'hB3D1, 16'hCCD4, 16'hCCD4, 16'hBC52, 16'hDD56, 16'hD516, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC515, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hC4D4, 16'hC4D5, 16'hBC93, 16'h9B4E, 16'hABD0, 16'hB451, 16'hD556, 16'hA410, 16'h7208, 16'hD4D3, 16'hD493, 16'hCC92, 16'hD493, 16'hC451, 16'h7A48, 16'h7248, 16'hCCD3, 16'h9B4D, 16'h930B, 16'h934D, 16'hABCF, 16'h7A8A, 16'hC556, 16'hC556, 16'hC516, 16'hC516, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hCD57, 16'hCD97, 16'hC556, 16'hCD97, 16'hCD97, 16'h9C51, 16'h72CB, 16'h834D, 16'hCE18, 16'hFFDF, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF6DB, 16'hD452, 16'hFE9B, 16'hFF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hFF5D, 16'hF6DB, 16'hF69B, 16'hF69B, 16'hDD97, 16'hC492, 16'hEE1A, 16'hFE9B, 16'hEE5A,
        16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE598, 16'hDD16, 16'hE597, 16'hEE5A, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF1D, 16'hED98, 16'hEDD9, 16'hFE9C, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE9C, 16'hF65B, 16'hF65B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE9B, 16'hED98, 16'hE516, 16'hFE5B, 16'hFE1A, 16'hFE1B, 16'hF65A, 16'hF65B, 16'hF65B, 16'hFE1A, 16'hF61A, 16'hFE1A, 16'hF61A, 16'hFE1B, 16'hDC94, 16'hED98, 16'hF61A, 16'hF5D9, 16'hF61A, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hEDD9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hBBD1, 16'hDD57, 16'hE5D9, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE5D8, 16'hFF5E, 16'hFF9F, 16'hF75D, 16'hFF5E, 16'hE619, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD97, 16'hDD97, 16'hDD97, 16'hCD15, 16'hCD15, 16'hDD97, 16'hC493, 16'hB412, 16'hDD56, 16'hB411, 16'hCD15, 16'hD556, 16'hCD15, 16'hCD15, 16'hCD15,
        16'hC515, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hC4D4, 16'hCCD5, 16'h9B4E, 16'hB411, 16'h9B4D, 16'hCD14, 16'hA3D0, 16'h828A, 16'hABD0, 16'hC492, 16'hD514, 16'hD4D3, 16'hD4D3, 16'h7A89, 16'h7A8A, 16'hCCD3, 16'h930C, 16'h8B0B, 16'h934D, 16'hABCF, 16'h7249, 16'hC515, 16'hC516, 16'hC515, 16'hC515, 16'hC516, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC596, 16'hBD55, 16'h9410, 16'h838D, 16'hACD3, 16'hD659, 16'hDE59, 16'hA451, 16'h9C0F, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD4D3, 16'hE597, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hFF5D, 16'hFF1D, 16'hF69B, 16'hF69B, 16'hFE9C, 16'hDD96, 16'hD596, 16'hF6DC, 16'hF69B, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hCCD5, 16'hED97, 16'hE598, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF1D, 16'hF69B, 16'hE516, 16'hFE9C, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hED56, 16'hED98, 16'hFE5B, 16'hF61A, 16'hF61A, 16'hF65B, 16'hFF9E, 16'hF69C, 16'hF69B, 16'hF69C, 16'hF61A, 16'hFE1A, 16'hFE1A, 16'hDC94, 16'hED98, 16'hF61A,
        16'hF61A, 16'hF5DA, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hEDD9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hAB4E, 16'hD515, 16'hE5D9, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE65A, 16'hF69C, 16'hE619, 16'hE619, 16'hE5D8, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD97, 16'hDD97, 16'hDD57, 16'hD556, 16'hCCD5, 16'hDD57, 16'hD556, 16'hB411, 16'hD516, 16'hC493, 16'hBC53, 16'hD556, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC515, 16'hC515, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hC4D4, 16'hCD15, 16'hB411, 16'hA38E, 16'h930D, 16'hB411, 16'hB451, 16'h61C6, 16'h82CB, 16'h5145, 16'hAB8F, 16'hD4D4, 16'hD4D4, 16'h7249, 16'h82CB, 16'hC492, 16'h930C, 16'h7207, 16'hABCF, 16'hABCF, 16'h7249, 16'hC515, 16'hBD16, 16'hC515, 16'hC515, 16'hC515, 16'hC516, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hBD15, 16'h838E, 16'h838E, 16'hBD54, 16'hBD55, 16'h9C51, 16'h93CF,
        16'hB514, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE618, 16'hCC53, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF5D,
        16'hFF1D, 16'hFF1D, 16'hFEDC, 16'hF69B, 16'hF6DD, 16'hF6DC, 16'hEE9A, 16'hFEDC, 16'hF6DC, 16'hF6DC, 16'hF69B, 16'hE5D8, 16'hE5D9, 16'hF65B, 16'hDD97, 16'hDD16, 16'hE557, 16'hF6DC, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFEDD, 16'hED97, 16'hED98, 16'hFE9C, 16'hFE1A, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hF61A, 16'hE515, 16'hF61A, 16'hFE1A, 16'hF61A, 16'hF61A, 16'hFEDC, 16'hFFDF, 16'hF65B, 16'hFF1D, 16'hFF9E, 16'hF65B, 16'hFE1A, 16'hFE1B, 16'hDC94, 16'hED98, 16'hF65B, 16'hF65C, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF61A, 16'hEDD9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D9, 16'hA34E, 16'hCCD4, 16'hE5D9, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hDD98, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hDD98, 16'hE598, 16'hDD98, 16'hDD97, 16'hDD97, 16'hDD57,
        16'hDD57, 16'hCD15, 16'hD515, 16'hD556, 16'hBC52, 16'hBC93, 16'hD515, 16'hABD0, 16'hCCD5, 16'hCD15, 16'hCD15, 16'hC515, 16'hC515, 16'hC515, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hC515, 16'hC4D4, 16'h9B4D, 16'h9B4E, 16'h9B8E, 16'hBC93, 16'h48C2, 16'hAC10, 16'hAC10, 16'h4080, 16'h9B8E, 16'hDD55, 16'h8ACB, 16'h7A49, 16'hC492, 16'h8ACB, 16'h7207, 16'hBC52, 16'h82CB, 16'h938E, 16'hCD56, 16'hBD15, 16'hBD16, 16'hC515, 16'hC515, 16'hBD16, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hAC93, 16'h834D, 16'h9C51, 16'hB514, 16'h9C50, 16'h6248, 16'h940F, 16'hF79D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5D, 16'hD493, 16'hF69B, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5D, 16'hFF9E, 16'hFFDF, 16'hF6DC, 16'hF6DC, 16'hFEDC, 16'hF69B, 16'hDDD8, 16'hD556, 16'hD556, 16'hEE5A, 16'hF69B, 16'hD515, 16'hE557, 16'hE5D8, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFEDD, 16'hF65B, 16'hE515, 16'hF65A, 16'hF61A, 16'hF61A, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5B, 16'hFE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hFE5B, 16'hED98, 16'hDCD5, 16'hFE5B, 16'hF61A, 16'hF61A,
        16'hF61A, 16'hF69C, 16'hFF5E, 16'hF65A, 16'hFF1D, 16'hFF9E, 16'hF65B, 16'hF61A, 16'hFE5B, 16'hDCD5, 16'hED98, 16'hF65B, 16'hF65B, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF61A, 16'hEE19, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hEDD9, 16'hAB4E, 16'hC452, 16'hEDD9, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hDD98, 16'hDD98, 16'hDD97, 16'hDD97, 16'hDD57, 16'hDD57, 16'hD516, 16'hCCD5, 16'hD556, 16'hC4D4, 16'hAB8F, 16'hCD16, 16'hB3D1, 16'hBC52, 16'hCD15, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hC4D4, 16'hCD15, 16'hABD0, 16'h9B8E, 16'h934D, 16'hC4D4, 16'h7A8A, 16'h7289, 16'hD514, 16'hA3CF, 16'h4080, 16'hB450, 16'h8ACB, 16'h7249, 16'hBC51, 16'h8289, 16'h7248, 16'hABCF, 16'h6A07, 16'hB492, 16'hC556, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD16,
        16'hC556, 16'hBD56, 16'hC556, 16'hB4D4, 16'h8B8F, 16'h9410, 16'hA492, 16'hACD3, 16'h940F, 16'h834C, 16'h838C, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hE5D7, 16'hDD56, 16'hFF5E, 16'hFF5E, 16'hFF5D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5D, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hFF9E, 16'hF6DC, 16'hEE5A, 16'hDD97, 16'hCD55, 16'hCD97, 16'hEE5A, 16'hFEDC, 16'hFEDC, 16'hE597, 16'hDD56, 16'hE597, 16'hF71D, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF1E, 16'hFEDD, 16'hED97, 16'hED97, 16'hF61A, 16'hEDD9, 16'hF61A, 16'hF61A, 16'hF65A, 16'hFE5B, 16'hFE5B, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hFE5B, 16'hE556, 16'hE556, 16'hFE1A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF65A, 16'hF619, 16'hFEDD, 16'hFF5D, 16'hF65A, 16'hF61A, 16'hFE5B, 16'hDCD5, 16'hED98, 16'hF61A, 16'hF61A, 16'hF5DA, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hEDD9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hEDD9, 16'hAB4E, 16'hB3D0, 16'hEDD9, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE598,
        16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hDD98, 16'hDD98, 16'hDD97, 16'hDD97, 16'hDD97, 16'hCD15, 16'hD516, 16'hD516, 16'hC4D4, 16'hD516, 16'hD556, 16'hABD0, 16'hC494, 16'hC493, 16'hA38F, 16'hCD15, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D5, 16'hC4D4, 16'hCD15, 16'hC493, 16'h934D, 16'h930D, 16'hB451, 16'hBC52, 16'h4000, 16'hB450, 16'hDD15, 16'h9B8E, 16'h61C6, 16'h7248, 16'h7249, 16'hB40F, 16'h69C6, 16'h8B0B, 16'h9B4D, 16'h7249, 16'hC515, 16'hC516, 16'hBD15, 16'hBD16, 16'hBD15, 16'hC515, 16'hBD16, 16'hBD16, 16'hBD56, 16'hAC92, 16'h834E, 16'hBD55, 16'hBD15, 16'h730D, 16'h9450, 16'hA4D2, 16'h93CF, 16'h5184, 16'hC596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'hCC93, 16'hF69B, 16'hFF1E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hEE5A, 16'hDD97, 16'hE5D8, 16'hEE9B, 16'hFEDC, 16'hF6DC, 16'hF6DC, 16'hF69B, 16'hCD15, 16'hE5D8, 16'hE619, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFEDD, 16'hF69B, 16'hD4D5, 16'hEDD8, 16'hE598, 16'hE598, 16'hE5D9, 16'hEDD9, 16'hEDD9, 16'hF61A,
        16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hFE1A, 16'hDCD4, 16'hF5D8, 16'hFE1A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF5DA, 16'hF619, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hFE1A, 16'hDCD5, 16'hED57, 16'hF61A, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hEDD9, 16'hEDD9, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hEDD9, 16'hABD0, 16'h8A8A, 16'hE5D8, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hDD98, 16'hDD98, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD97, 16'hD556, 16'hCCD4, 16'hD516, 16'hCCD5, 16'hCD15, 16'hD516, 16'hBC52, 16'hABD0, 16'hD515, 16'hA38F, 16'hC4D4, 16'hCD15, 16'hC4D5, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hCD15, 16'h934D, 16'h934D, 16'hAC10, 16'hCD15, 16'h934D, 16'h61C7, 16'hCCD4, 16'hD515, 16'h7289, 16'h4903, 16'h6A08,
        16'hA38D, 16'h61C6, 16'hA38E, 16'h69C6, 16'hAC51, 16'hC556, 16'hBD15, 16'hBD15, 16'hBD16, 16'hBD15, 16'hC515, 16'hBD16, 16'hBD16, 16'hC556, 16'hAC93, 16'h9410, 16'hB514, 16'hC556, 16'hBD55, 16'h6B0B, 16'h838E, 16'hC596, 16'h838D, 16'h7B4B, 16'hF79D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDD55, 16'hDD56, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFF5D, 16'hF6DC, 16'hDDD8, 16'hDD97, 16'hF69B, 16'hF6DD, 16'hF6DC, 16'hFEDC, 16'hDD97, 16'hDD97, 16'hDD97, 16'hF71D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF1E, 16'hFEDC, 16'hEDD8, 16'hDCD5, 16'hE598, 16'hDD57, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE5D8, 16'hEDD9, 16'hEDD9, 16'hF619, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF5D9, 16'hCC52, 16'hED98, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF619, 16'hF61A, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF619, 16'hF5D9, 16'hF61A, 16'hDCD5, 16'hE557, 16'hF61A, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE5D9, 16'hB3D1,
        16'h7104, 16'hDD56, 16'hE5D9, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hDD98, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD57, 16'hDD57, 16'hDD57, 16'hCCD5, 16'hCD15, 16'hCD15, 16'hCCD4, 16'hCD15, 16'hCCD4, 16'hA34E, 16'hCCD4, 16'hB411, 16'hB452, 16'hCD15, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hCD15, 16'hAC11, 16'h7249, 16'h934D, 16'hB492, 16'hC4D3, 16'h7208, 16'h82CB, 16'hD555, 16'hB451, 16'h2800, 16'h7289, 16'h7A48, 16'h6A48, 16'h828A, 16'h830C, 16'hC555, 16'hBD16, 16'hC515, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD16, 16'hBD16, 16'hBD16, 16'hC556, 16'hAC93, 16'h72CB, 16'h7B4D, 16'h9C52, 16'h6ACC, 16'h5249, 16'h9C51, 16'hA492, 16'h5181, 16'hD658, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'hC452, 16'hF69B, 16'hFF1E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5D, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hF6DC, 16'hE619, 16'hDDD8, 16'hF6DC, 16'hFF1D, 16'hF6DC, 16'hEE9B, 16'hEE5B, 16'hD556, 16'hE5D8, 16'hDDD7, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5E,
        16'hFF1E, 16'hFEDD, 16'hFE9C, 16'hDD56, 16'hDD56, 16'hE598, 16'hDD57, 16'hDD98, 16'hDD98, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hEDD8, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hE556, 16'hC410, 16'hDCD5, 16'hF5D9, 16'hF61A, 16'hF619, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hEDD9, 16'hEDD9, 16'hF5D9, 16'hEDD9, 16'hEDD9, 16'hF61A, 16'hD4D5, 16'hDD16, 16'hF61A, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE5D9, 16'hB3D1, 16'h81C7, 16'hC493, 16'hE5D9, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hDD98, 16'hDD98, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD57, 16'hD556, 16'hD556, 16'hDD56, 16'hD515, 16'hC494, 16'hCD15, 16'hC4D4, 16'hCCD5, 16'hCD15, 16'hABD0, 16'hBC52, 16'hC493, 16'hA3CF, 16'hCD15, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D5, 16'hC4D5, 16'hC4D5,
        16'hC515, 16'hBC93, 16'h61C7, 16'h6A49, 16'h728A, 16'h8B0C, 16'h8B0C, 16'h40C1, 16'h938D, 16'hBC92, 16'h4944, 16'h7289, 16'h6207, 16'h7207, 16'h7A49, 16'hBCD3, 16'hC556, 16'hBD15, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hBD16, 16'hBD16, 16'hBD16, 16'hBD56, 16'hB4D4, 16'h7B4D, 16'h4186, 16'h730C, 16'h83CF, 16'h6ACC, 16'h62CB, 16'hA4D3, 16'h6ACA, 16'hA491, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD596, 16'hD555, 16'hFF5D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hF6DB, 16'hD5D7, 16'hD596, 16'hF69B, 16'hF6DC, 16'hEE5A, 16'hD596, 16'hCD55, 16'hDDD8, 16'hDD96, 16'hDD56, 16'hDD56, 16'hEEDC, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5E, 16'hFF1E, 16'hFF1D, 16'hFEDC, 16'hF61A, 16'hCC93, 16'hDD57, 16'hDD57, 16'hDD97, 16'hDD97, 16'hDD98, 16'hDD97, 16'hDD97, 16'hDD97, 16'hE598, 16'hE598, 16'hE5D8, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hCC93, 16'hC411, 16'hD4D4, 16'hF5D9, 16'hEE1A, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hD4D5, 16'hD515, 16'hEDD9, 16'hE598, 16'hE598, 16'hE5D8, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598,
        16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hEDD9, 16'hB411, 16'h7986, 16'hB3D0, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hDD98, 16'hDD98, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD57, 16'hD556, 16'hD556, 16'hD516, 16'hD516, 16'hD516, 16'hC493, 16'hCCD4, 16'hC4D4, 16'hCCD4, 16'hCD15, 16'hBC52, 16'hABD0, 16'hCCD4, 16'hA38F, 16'hC4D4, 16'hCD15, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D5, 16'hC515, 16'hC4D4, 16'h828B, 16'h69C7, 16'h8B0C, 16'h7289, 16'h59C6, 16'h6207, 16'h4102, 16'h7A89, 16'h59C6, 16'h4944, 16'h5986, 16'h7A89, 16'hB451, 16'hCD56, 16'hC556, 16'hC556, 16'hBD14, 16'hB493, 16'hA411, 16'h9BD0, 16'hB514, 16'hC556, 16'hBD16, 16'hBD56, 16'hBD56, 16'hC556, 16'hA493, 16'h5208, 16'hACD3, 16'hC597, 16'hB555, 16'hBD56, 16'hC597, 16'h9410, 16'h6206, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hC452, 16'hEE5A, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5D, 16'hF71D, 16'hEE9A, 16'hD596, 16'hCD56, 16'hE619, 16'hF69B, 16'hE5D8, 16'hCD15, 16'hD597,
        16'hE5D8, 16'hF69B, 16'hF69B, 16'hC4D3, 16'hE5D8, 16'hDD56, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF1E, 16'hFF1D, 16'hFEDC, 16'hFE9C, 16'hDD56, 16'hCCD4, 16'hDD97, 16'hDD57, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD97, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hEDD9, 16'hBC11, 16'hCC51, 16'hD493, 16'hF619, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hE598, 16'hE5D9, 16'hD4D5, 16'hCCD4, 16'hDD98, 16'hDD57, 16'hDD57, 16'hDD97, 16'hDD97, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD97, 16'hE598, 16'hE598, 16'hE5D8, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hEDD9, 16'hC452, 16'h7185, 16'hA30D, 16'hDD97, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hDD98, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD57, 16'hD556, 16'hD516, 16'hCD15, 16'hCD15, 16'hCD15, 16'hD516, 16'hCCD4, 16'hC494, 16'hCCD4, 16'hC4D4, 16'hCCD5, 16'hC494, 16'hA34E,
        16'hC493, 16'hABD0, 16'hBC93, 16'hCD15, 16'hC4D5, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D4, 16'hCD15, 16'hAC10, 16'h6145, 16'h934C, 16'h934C, 16'h7A8A, 16'h5144, 16'h5144, 16'h4103, 16'h5185, 16'h6A48, 16'h59C6, 16'h4104, 16'h5A07, 16'h938E, 16'h938E, 16'h8B4D, 16'h7249, 16'h6A07, 16'h8ACA, 16'h8ACA, 16'h7289, 16'hACD4, 16'hC556, 16'hC556, 16'hBD56, 16'hBD56, 16'hBD55, 16'h6ACB, 16'h838E, 16'hB515, 16'hBD97, 16'hBD56, 16'hBD97, 16'hA493, 16'h59C6, 16'hC596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9B, 16'hCCD3, 16'hFEDC, 16'hFF1E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hE65A, 16'hDDD7, 16'hEE5A, 16'hF6DC, 16'hFEDC, 16'hE65A, 16'hDDD8, 16'hF69B, 16'hFEDC, 16'hF6DC, 16'hF6DC, 16'hE5D8, 16'hD596, 16'hDDD8, 16'hE619, 16'hFFDF, 16'hFF9F, 16'hFF5F, 16'hFF1E, 16'hFF1D, 16'hFEDC, 16'hF69B, 16'hF65A, 16'hC452, 16'hD516, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD97, 16'hDD97, 16'hE598, 16'hE598, 16'hE598, 16'hB3D0, 16'hC411, 16'hC452, 16'hF5D9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hE5D8, 16'hE598, 16'hE598,
        16'hE598, 16'hCCD5, 16'hCC94, 16'hDD57, 16'hD556, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hD556, 16'hD556, 16'hD556, 16'hDD57, 16'hDD57, 16'hDD98, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE5D8, 16'hC452, 16'h6945, 16'h9ACB, 16'hC4D4, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD57, 16'hD556, 16'hD516, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hC494, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hCCD4, 16'hABD0, 16'hBC52, 16'hBC52, 16'hB411, 16'hCD15, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D4, 16'hC515, 16'hC4D3, 16'h69C7, 16'h9B8F, 16'hCD14, 16'hC493, 16'hBC92, 16'hB451, 16'h8B0B, 16'h6207, 16'h59C6, 16'h6207, 16'h934C, 16'h82CA, 16'h4040, 16'h7A88, 16'h9B4C, 16'hABCF, 16'hCC92, 16'hD4D3, 16'hD493, 16'hAB8E, 16'h51C6, 16'hAC93, 16'hC556, 16'hBD56, 16'hBD56, 16'hC557, 16'h9C11, 16'h28C1, 16'h730C,
        16'hA4D3, 16'hBD56, 16'hBD56, 16'hB555, 16'h6249, 16'h8BCE, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDDD8, 16'hCCD3, 16'hFEDD,
        16'hFF1D, 16'hFF1C, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hF6DC, 16'hF69B, 16'hF69B, 16'hF69C, 16'hFEDC, 16'hF69C, 16'hF69B, 16'hF69B, 16'hF69B, 16'hCD14, 16'hE619, 16'hCD15, 16'hF71D, 16'hFF9F, 16'hFF5F, 16'hFF1E, 16'hFF1E, 16'hFEDD, 16'hFEDC, 16'hF65B, 16'hE597, 16'hC452, 16'hD557, 16'hD557, 16'hD557, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hD516, 16'hD557, 16'hDD57, 16'hDD57, 16'hE598, 16'hE557, 16'hAB4E, 16'hB38F, 16'hC493, 16'hEDD9, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hDD97, 16'hDD98, 16'hD4D5, 16'hC493, 16'hD557, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD516, 16'hD516, 16'hD556, 16'hD556, 16'hD556, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD97, 16'hDD97, 16'hDD97, 16'hE598, 16'hC493, 16'h5842, 16'h9B0C, 16'hB411, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hE598, 16'hDD98, 16'hDD98, 16'hE598, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD57, 16'hDD57, 16'hD556, 16'hCD16,
        16'hCD15, 16'hCCD5, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hCCD5, 16'hC494, 16'hC494, 16'hC4D4, 16'hC4D4, 16'hCCD4, 16'hB411, 16'hABD0, 16'hC493, 16'hA3CF, 16'hCD15, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D4, 16'hCD15, 16'h8B0C, 16'h8B0D, 16'hCD56, 16'hCD15, 16'hCD56, 16'hBCD3, 16'h7A89, 16'h5185, 16'h3882, 16'h5185, 16'h6A08, 16'h8ACA, 16'h7248, 16'h5185, 16'h934C, 16'hA38E, 16'hBC10, 16'hBC51, 16'hC451, 16'hCC92, 16'h9B8D, 16'h7B4D, 16'hC556, 16'hC556, 16'hC556, 16'hC557, 16'hACD4, 16'h628A, 16'h7B4D, 16'h838F, 16'hBD56, 16'hB556, 16'hBD56, 16'h8BCF, 16'h5182, 16'hDE99, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hD555, 16'hC452, 16'hF69B, 16'hF6DC, 16'hF6DC, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69C, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hEE9B, 16'hEE19, 16'hCD15, 16'hE619, 16'hD556, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF1E, 16'hFF1D, 16'hFEDC, 16'hFE9B, 16'hF61A, 16'hCCD5, 16'hC4D4, 16'hD557, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD15, 16'hD556, 16'hDD57, 16'hDD57, 16'hE597, 16'hD4D5, 16'hA30D, 16'hB3D0,
        16'hCC94, 16'hE598, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD57, 16'hDD97, 16'hE598, 16'hDD97, 16'hDD97, 16'hDD57, 16'hDD57, 16'hDD57, 16'hCCD4, 16'hC493, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'hD556, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hE598, 16'hC493, 16'h79C8, 16'h9ACC, 16'hAB4E, 16'hDD97, 16'hE598, 16'hDD98, 16'hE598, 16'hDD97, 16'hDD97, 16'hDD57, 16'hDD57, 16'hDD57, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD557, 16'hD556, 16'hCD15, 16'hCCD5, 16'hCCD5, 16'hCCD5, 16'hCCD5, 16'hCCD5, 16'hCCD5, 16'hCCD4, 16'hC493, 16'hC494, 16'hC494, 16'hC4D4, 16'hC452, 16'hA38E, 16'hC4D4, 16'hA38F, 16'hC4D4, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D4, 16'hCD15, 16'hA3D0, 16'h7249, 16'hC515, 16'hCD56, 16'hB452, 16'h5985, 16'h7248, 16'h59C6, 16'h5185, 16'h5145, 16'h4944, 16'h38C1, 16'h7248, 16'h6207, 16'h28C2, 16'h72CB, 16'h7289,
        16'h7289, 16'h7248, 16'h7A8A, 16'h830B, 16'h51C6, 16'h72CC, 16'h9C11, 16'hB515, 16'hC596, 16'hC556, 16'h834E, 16'h9C51, 16'hBD56, 16'hB515, 16'hB515, 16'hBD56, 16'hA492, 16'h48C0, 16'hBD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hCD14, 16'hD515, 16'hFEDC, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hD596, 16'hDDD7, 16'hDD56, 16'hEE5A, 16'hFFDF, 16'hFF5F, 16'hFF1E, 16'hFF1D, 16'hFEDD, 16'hFE9C, 16'hF65A, 16'hE598, 16'hC493, 16'hCD15, 16'hD557, 16'hD516, 16'hD556, 16'hD556, 16'hD516, 16'hD516, 16'hD556, 16'hD556, 16'hCD15, 16'hCCD5, 16'hD516, 16'hD516, 16'hD556, 16'hDD57, 16'hC453, 16'hA34E, 16'hA34E, 16'hCC94, 16'hDD57, 16'hD556, 16'hD556, 16'hD556, 16'hD516, 16'hD516, 16'hD556, 16'hD556, 16'hD556, 16'hD516, 16'hD516, 16'hD556, 16'hCCD4, 16'hC494, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hCD15, 16'hD516, 16'hD516, 16'hD556, 16'hD556, 16'hDD57, 16'hDD57, 16'hDD57, 16'hC493, 16'h8ACB, 16'hA34D, 16'h9A8B, 16'hCCD4, 16'hE598, 16'hDD97, 16'hDD97, 16'hDD57,
        16'hDD57, 16'hD556, 16'hD556, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'hD516, 16'hD556, 16'hD556, 16'hCD15, 16'hCCD5, 16'hCCD5, 16'hCCD5, 16'hCCD5, 16'hCCD5, 16'hCCD4, 16'hCCD4, 16'hC493, 16'hC493, 16'hC494, 16'hC4D4, 16'hC493, 16'h9B4E, 16'hC493, 16'hABD0, 16'hBC93, 16'hC515, 16'hC4D4, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D4, 16'hCD15, 16'hBC93, 16'h61C7, 16'hBCD3, 16'hAC51, 16'h50C1, 16'h9B4C, 16'h828A, 16'h7A49, 16'h6A07, 16'h6A48, 16'h59C6, 16'h6A48, 16'h6A07, 16'hA38D, 16'h6A07, 16'h93CF, 16'hBCD4, 16'hAC93, 16'hA412, 16'hA452, 16'h9BD0, 16'h7A8B, 16'h40C3, 16'h72CB, 16'h72CC, 16'h9C11, 16'hB4D4, 16'h9C51, 16'h5A49, 16'hB4D5, 16'hB516, 16'hB515, 16'hBD56, 16'hACD3, 16'h72CA, 16'h8B8D, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF6DC, 16'hBC11, 16'hDD97, 16'hF69C, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hCD14, 16'hE619, 16'hCCD4, 16'hFF1D, 16'hFF9F, 16'hFF5E, 16'hFF1D, 16'hFEDC, 16'hFEDC, 16'hF69B, 16'hEE19, 16'hD516, 16'hC452, 16'hD516, 16'hCD16, 16'hD516, 16'hD516, 16'hD516, 16'hD516,
        16'hD516, 16'hD516, 16'hD556, 16'hCCD5, 16'hCD15, 16'hD516, 16'hD516, 16'hD556, 16'hDD57, 16'hABD0, 16'hAB8E, 16'hA34D, 16'hC493, 16'hDD57, 16'hD556, 16'hD556, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hCD15, 16'hD516, 16'hCCD5, 16'hC493, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'hD516, 16'hCD15, 16'hD515, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'hD556, 16'hDD57, 16'hC494, 16'hA34D, 16'hC451, 16'h8A09, 16'hBC11, 16'hDD97, 16'hDD57, 16'hDD57, 16'hDD57, 16'hD556, 16'hD556, 16'hD516, 16'hD556, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'hCCD5, 16'hCCD4, 16'hD556, 16'hCD15, 16'hCCD5, 16'hCCD5, 16'hCCD4, 16'hCCD5, 16'hCCD5, 16'hCCD5, 16'hCCD4, 16'hC494, 16'hC493, 16'hC494, 16'hC494, 16'hCCD4, 16'hABD0, 16'hB411, 16'hBC52, 16'hB451, 16'hCD15, 16'hC4D4, 16'hC515, 16'hC4D5, 16'hC4D5, 16'hC515, 16'hC515, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hC4D4, 16'h7ACB, 16'h7ACA, 16'h5145, 16'hA38D,
        16'hABCE, 16'h69C7, 16'h9B4C, 16'h61C6, 16'h82CB, 16'h5185, 16'h7289, 16'h59C6, 16'hA38D, 16'h9B4C, 16'h4103, 16'hA451, 16'hC516, 16'hBCD5, 16'hBCD4, 16'hBCD5, 16'h9B8F, 16'h6186, 16'h9C10, 16'hAC93, 16'h93D0, 16'h838E, 16'h7B4D, 16'h7B4D, 16'hACD4, 16'hB515, 16'hB515, 16'hBD56, 16'hB515, 16'h834E, 16'h7ACA, 16'hD618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hCD55, 16'hC493, 16'hBC51, 16'hB411, 16'hE5D8, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hE618, 16'hD556, 16'hE5D8, 16'hD556, 16'hFF5F, 16'hFF5E, 16'hFF1E, 16'hFEDC, 16'hFEDC, 16'hFE9C, 16'hF65A, 16'hE5D8, 16'hCCD5, 16'hBC52, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hCD15, 16'hC494, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hDD57, 16'hA34E, 16'hABCF, 16'hAB8E, 16'hCCD4, 16'hD556, 16'hD556, 16'hD556, 16'hD516, 16'hCD15, 16'hD516, 16'hCD15, 16'hCD15, 16'hD516, 16'hD516, 16'hCD15, 16'hD516, 16'hCCD5, 16'hC493, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'hD516, 16'hCD15, 16'hCD15, 16'hD516, 16'hD516, 16'hD516,
        16'hD516, 16'hD516, 16'hDD56, 16'hCCD4, 16'h9B0C, 16'hC493, 16'h9B0C, 16'hAB8E, 16'hDD56, 16'hDD57, 16'hD556, 16'hD556, 16'hD556, 16'hD516, 16'hD516, 16'hD556, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hCD15, 16'hC493, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD5, 16'hCCD5, 16'hCCD4, 16'hC4D4, 16'hC493, 16'hC493, 16'hC494, 16'hC4D4, 16'hB452, 16'hA38F, 16'hBC52, 16'hA3D0, 16'hC515, 16'hC4D4, 16'hC515, 16'hC4D5, 16'hC4D5, 16'hC515, 16'hC515, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hCD15, 16'h934E, 16'h3800, 16'hA38D, 16'hC490, 16'h5945, 16'hA34D, 16'hAB8E, 16'h5186, 16'hA38E, 16'h61C6, 16'h7249, 16'h59C6, 16'h9B8D, 16'hC491, 16'h5985, 16'h6207, 16'h9BD0, 16'hBD15, 16'hBCD4, 16'hB494, 16'h8B0D, 16'h8B0C, 16'h9BD0, 16'hBD16, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hB515, 16'hB515, 16'hBD15, 16'hBD15, 16'hBD56, 16'h93D0, 16'h830C, 16'hAC92, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hCD15, 16'hA2CC, 16'hC452, 16'hEE19, 16'hEE5A, 16'hDD97, 16'hEE5A, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hD555, 16'hE619, 16'hCD14, 16'hE659, 16'hFF9F, 16'hFF5E, 16'hFF1D, 16'hF69C,
        16'hF69B, 16'hF65B, 16'hEE19, 16'hDD97, 16'hBC52, 16'hC4D4, 16'hD556, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hD516, 16'hD516, 16'hC4D5, 16'hC4D4, 16'hD516, 16'hD516, 16'hD516, 16'hCD15, 16'hDD56, 16'h9B4E, 16'hBC11, 16'hA38E, 16'hCCD5, 16'hD556, 16'hD556, 16'hD516, 16'hD516, 16'hCD15, 16'hD516, 16'hCD15, 16'hCD15, 16'hD516, 16'hD516, 16'hCD15, 16'hD516, 16'hCCD5, 16'hC493, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD516, 16'hCD15, 16'hCD15, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'hD4D5, 16'h92CB, 16'hD515, 16'h92CC, 16'h9ACB, 16'hD4D4, 16'hDD97, 16'hD556, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hBC52, 16'hC4D4, 16'hCD16, 16'hCCD5, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hC494, 16'hC493, 16'hC493, 16'hC493, 16'hC494, 16'hC493, 16'h9B4E, 16'hBC52, 16'hA3D0, 16'hC4D5, 16'hC515, 16'hC515, 16'hC515,
        16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D4, 16'hCD15, 16'hA3D0, 16'h61C6, 16'hCC91, 16'h7A48, 16'h7208, 16'hC451, 16'h930B, 16'h3944, 16'hAC0F, 16'h8ACA, 16'h7248, 16'h4944, 16'h6A07, 16'hCD12, 16'h82CA, 16'h7248, 16'h82CA, 16'h938E, 16'hBCD4, 16'hAC93, 16'h6A49, 16'h828A, 16'h938F, 16'hBD15, 16'hB4D4, 16'hBD15, 16'hBD15, 16'hB4D5, 16'hB515, 16'hB515, 16'hBD15, 16'hBD15, 16'hBD56, 16'hA452, 16'h830C, 16'hA40F, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hD515, 16'hCC93, 16'hEE1A, 16'hFE9B, 16'hEE5B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF65A, 16'hD555, 16'hE619, 16'hC493, 16'hFF1D, 16'hFF5E, 16'hFF1D, 16'hF6DC, 16'hF69B, 16'hF69B, 16'hF65A, 16'hE5D9, 16'hD515, 16'hBC52, 16'hCD15, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hC494, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hD516, 16'hC4D4, 16'h61C7, 16'hBC51, 16'h9B4D, 16'hCCD5, 16'hD556, 16'hD556, 16'hD516, 16'hD516, 16'hCD15, 16'hD516, 16'hCD15, 16'hCD15, 16'hD516, 16'hD516, 16'hCD15, 16'hD516, 16'hD515, 16'hC453, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556,
        16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD516, 16'hCD15, 16'hCD15, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'hCCD5, 16'h8208, 16'hEDD8, 16'hB411, 16'h9248, 16'hBC11, 16'hDD97, 16'hD556, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'hC4D4, 16'hBC53, 16'hCD15, 16'hCCD5, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hCCD4, 16'hC4D4, 16'hC494, 16'hC493, 16'hBC53, 16'hC493, 16'hC493, 16'hCCD4, 16'h9B4E, 16'hB451, 16'hABD0, 16'hC4D4, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D4, 16'hC515, 16'hB452, 16'h7208, 16'h7248, 16'h5104, 16'hB410, 16'hCC92, 16'h7A8A, 16'h1881, 16'hB450, 16'h930C, 16'h82CB, 16'h51C6, 16'h38C1, 16'hBC51, 16'hBC91, 16'h5101, 16'hB40F, 16'h9B4E, 16'h6A49, 16'h830C, 16'h7A8A, 16'h828A, 16'h93CF, 16'hBD15, 16'hB514, 16'hBD15, 16'hBD15, 16'hB515, 16'hB515, 16'hB515, 16'hB515, 16'hBD15, 16'hBD56, 16'hB4D4, 16'h830C, 16'hA3CF,
        16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hE5D7, 16'hBC10, 16'hD515, 16'hEE19, 16'hF69B, 16'hF69B, 16'hF69C, 16'hEE9B,
        16'hF69B, 16'hEE9B, 16'hF6DC, 16'hE618, 16'hD556, 16'hDD97, 16'hCD15, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hF69B, 16'hF65B, 16'hF65A, 16'hEE19, 16'hE598, 16'hCCD4, 16'hB452, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD16, 16'hCCD5, 16'hC493, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hD556, 16'hABD0, 16'h48C2, 16'hBC92, 16'h930C, 16'hCD15, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hCD15, 16'hD516, 16'hCD15, 16'hCD15, 16'hCD15, 16'hD516, 16'hCD15, 16'hCD16, 16'hCD15, 16'hC453, 16'hD516, 16'hD556, 16'hD556, 16'hD556, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hCD15, 16'hCD15, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'hD515, 16'h8208, 16'hE597, 16'hD515, 16'h8A08, 16'hA34E, 16'hD556, 16'hDD57, 16'hD516, 16'hD516, 16'hD556, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hCD15, 16'hBC52, 16'hCD15, 16'hCCD5, 16'hCCD4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC494,
        16'hC494, 16'hBC52, 16'hC493, 16'hC493, 16'hCCD4, 16'hA38F, 16'hB411, 16'hB411, 16'hBC93, 16'hC515, 16'hC514, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hC515, 16'hC4D4, 16'h6A08, 16'h4904, 16'hABCF, 16'hCCD3, 16'hC451, 16'h51C6, 16'h4145, 16'hA3CE, 16'hA38E, 16'h938D, 16'h7ACB, 16'h6207, 16'h61C7, 16'hBC50, 16'h7247, 16'h9B4D, 16'hD4D4, 16'h9B8E, 16'h61C7, 16'hAC10, 16'h7A8A, 16'hA411, 16'hBD15, 16'hB4D5, 16'hB515, 16'hBD15, 16'hB515, 16'hB515, 16'hB514, 16'hB515, 16'hB515, 16'hBD15, 16'hBD56, 16'h8B8E, 16'h938D, 16'hC555, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hCD15, 16'hC493, 16'hD556, 16'hEE19, 16'hEE5A, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF69B, 16'hD555, 16'hEE59, 16'hCC93, 16'hE619, 16'hFF5E, 16'hFF1D, 16'hF6DC, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hE5D9, 16'hDD97, 16'hBC53, 16'hBC93, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD16, 16'hC494, 16'hC4D4, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hD515, 16'h9B4D, 16'h7A08, 16'hBC92, 16'h9B4D, 16'hCD15, 16'hD516, 16'hD516, 16'hD516, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15,
        16'hCD15, 16'hD516, 16'hD516, 16'hCD15, 16'hCD15, 16'hCD16, 16'hC453, 16'hCD16, 16'hD556, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hCD15, 16'hCD15, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'h92CB, 16'hDD56, 16'hF61A, 16'h9B0C, 16'h8A49, 16'hCCD4, 16'hDD97, 16'hD516, 16'hD516, 16'hD556, 16'hD556, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hCD15, 16'hD516, 16'hBC53, 16'hC494, 16'hCD15, 16'hCCD4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC494, 16'hC494, 16'hC453, 16'hBC52, 16'hC493, 16'hC494, 16'hB411, 16'hABCF, 16'hB411, 16'hB411, 16'hCD15, 16'hC4D4, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hCCD5, 16'h82CB, 16'h7A8A, 16'hCCD3, 16'hD4D3, 16'h9B4D, 16'h000, 16'h7B0B, 16'h934D, 16'hA3CF, 16'h8B4D, 16'h8B4D, 16'h8B4C, 16'h728A, 16'h48C3, 16'h82CA, 16'h6A07, 16'hBC50, 16'hCCD4, 16'hCCD4, 16'hBC51, 16'h6A07, 16'hB493, 16'hBD15,
        16'hB4D5, 16'hBD15, 16'hBD15, 16'hB515, 16'hB515, 16'hB515, 16'hB515, 16'hBD15, 16'hBD15, 16'hBD56, 16'h9C10, 16'h8B4D, 16'hB492, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hE5D8, 16'hCC93, 16'hC452, 16'hD556, 16'hE5D8, 16'hEE5A, 16'hF69B, 16'hEE5A, 16'hD555, 16'hEE5A, 16'hC492, 16'hF69B, 16'hFF5E, 16'hFF1D, 16'hF69C, 16'hEE1A, 16'hEE1A, 16'hE5D9, 16'hE5D8, 16'hDD57, 16'hB411, 16'hC4D4, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC494, 16'hCCD5, 16'hCD15, 16'hCD15, 16'hCD15, 16'hD516, 16'hBC92, 16'h92CB, 16'hA34D, 16'hBC92, 16'h9B8E, 16'hCD15, 16'hD516, 16'hD516, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hD516, 16'hD516, 16'hCD15, 16'hCD15, 16'hD516, 16'hC493, 16'hCD15, 16'hD556, 16'hD516, 16'hD516, 16'hCD16, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hCD15, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hDD56, 16'h9B0C, 16'hCCD3, 16'hFE9B, 16'hBC51, 16'h81C7, 16'hABD0, 16'hDD97, 16'hD516, 16'hCD15, 16'hD556, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516,
        16'hCD15, 16'hD516, 16'hCCD4, 16'hBC53, 16'hCD15, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC494, 16'hC494, 16'hC493, 16'hB411, 16'hC493, 16'hC493, 16'hBC52, 16'hA38E, 16'hBC11, 16'hAC11, 16'hCD15, 16'hC4D4, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D5, 16'hCD15, 16'h938E, 16'h7208, 16'hCC93, 16'hABCF, 16'h5186, 16'h4945, 16'h8B4C, 16'hA40F, 16'hA410, 16'h934D, 16'hA3CF, 16'h82CB, 16'hCCD3, 16'h934C, 16'h59C6, 16'h51C6, 16'h5984, 16'h8B0B, 16'hC493, 16'hA38E, 16'h6A07, 16'hB4D4, 16'hBD15, 16'hB514, 16'hB514, 16'hBD14, 16'hBD15, 16'hBD15, 16'hBD14, 16'hB4D4, 16'hB515, 16'hBD15, 16'hBD56, 16'hA492, 16'h834D, 16'hB491, 16'hDE99, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hE69B, 16'hDE59, 16'hCD96, 16'hCD15, 16'hCD14, 16'hCCD4, 16'hCD15, 16'hDD97, 16'hBC51, 16'hB451, 16'hEE19, 16'hF69B, 16'hE619, 16'hD555, 16'hE597, 16'hCCD4, 16'hFF1D, 16'hFF1D, 16'hFEDD, 16'hEE5B, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hDD98, 16'hD516, 16'hB411, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hC493, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hD556, 16'h9B8F,
        16'hABCF, 16'hA38E, 16'hB410, 16'h930C, 16'hCD15, 16'hD516, 16'hD516, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD16, 16'hCD15, 16'hCD15, 16'hD516, 16'hD516, 16'hCD15, 16'hCD15, 16'hD556, 16'hC493, 16'hCCD5, 16'hD516, 16'hD516, 16'hD516, 16'hCD16, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hCD15, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hDD56, 16'hA34D, 16'hBC51, 16'hFE9B, 16'hDD56, 16'h8A08, 16'h930B, 16'hCD15, 16'hD556, 16'hCD15, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hC493, 16'hCCD4, 16'hC4D4, 16'hCCD4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC493, 16'hC493, 16'hBC52, 16'hBC52, 16'hC493, 16'hC493, 16'h9B0D, 16'hB410, 16'hABD0, 16'hC515, 16'hC514, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D5, 16'hCD15, 16'hAC11, 16'h5144, 16'h930C, 16'h69C7, 16'h6A48, 16'h7A8A, 16'h8B4C, 16'hA410, 16'hA410, 16'h934E, 16'hAC10,
        16'h82CB, 16'hA3CF, 16'hD554, 16'hBC91, 16'h5186, 16'h82CB, 16'h6A08, 16'h6A06, 16'h61C6, 16'h9BCF, 16'hBD15, 16'hB4D4, 16'hB514, 16'hB514, 16'hB514, 16'hBD14, 16'hBD15, 16'hBD14, 16'hB4D4, 16'hB515, 16'hBD15, 16'hBD56, 16'hB4D4, 16'h72CA, 16'hC554, 16'hCDD6, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hC4D4, 16'hC4D4, 16'hD515, 16'hDD56, 16'hE618, 16'hFF1D, 16'hFF1D, 16'hCD15, 16'hC492, 16'hEE19, 16'hEE5A, 16'hF69B, 16'hDD96, 16'hE5D8, 16'hCD15, 16'hCD15, 16'hFF5E, 16'hFF1D, 16'hFEDC, 16'hEE1A, 16'hE5D9, 16'hE5D8, 16'hDD98, 16'hDD97, 16'hCCD4, 16'hB411, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC4D4, 16'hC4D4, 16'hCD15, 16'hCCD5, 16'hCD15, 16'hCD15, 16'hD555, 16'h930C, 16'hC492, 16'h8ACB, 16'hBC51, 16'h934D, 16'hCD15, 16'hD516, 16'hD516, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hD516, 16'hCD15, 16'hCD15, 16'hD556, 16'hC493, 16'hC4D4, 16'hD556, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hCD15, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hDD56, 16'hAB8F, 16'hB410, 16'hFE9C, 16'hF65A,
        16'h9B0B, 16'h8248, 16'hB451, 16'hDD56, 16'hCD15, 16'hCD15, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC493, 16'hC4D4, 16'hCCD4, 16'hC4D4, 16'hC4D4, 16'hC494, 16'hC494, 16'hC494, 16'hC4D4, 16'hC4D4, 16'hC494, 16'hBC93, 16'hB411, 16'hC493, 16'hCC93, 16'h9B4E, 16'hB3D0, 16'hABD0, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D4, 16'hC515, 16'hBC93, 16'h5986, 16'h51C6, 16'h9BCE, 16'h9B8D, 16'h7248, 16'h938E, 16'hA410, 16'h9BCF, 16'h9BCF, 16'h9B8F, 16'hAC11, 16'h7A49, 16'hC492, 16'hD514, 16'h9B8D, 16'h830C, 16'hBD14, 16'hB493, 16'hB4D3, 16'hBD14, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'hB514, 16'hBD15, 16'hBD15, 16'hB4D4, 16'hB515, 16'hBD15, 16'hBD15, 16'hBD55, 16'h728A, 16'hBD55, 16'hD5D7, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hE659, 16'hD5D7, 16'hDE18, 16'hE61A, 16'hABD0, 16'hCCD4, 16'hEE19, 16'hF65A, 16'hF69B, 16'hEE5A, 16'hCCD4, 16'hF69B, 16'hC493, 16'hE619, 16'hFF5E, 16'hFF1D, 16'hF69C, 16'hE5D9, 16'hE5D8, 16'hDD98, 16'hDD97, 16'hDD97, 16'hBC52, 16'hBC52, 16'hCD15, 16'hCCD5, 16'hCD15, 16'hCD15,
        16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC494, 16'hCCD5, 16'hCCD5, 16'hCCD5, 16'hCD15, 16'hCD16, 16'hC4D3, 16'h9B0D, 16'hDD56, 16'h92CB, 16'hC492, 16'h8B0C, 16'hCD15, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hD556, 16'hC494, 16'hC494, 16'hD556, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hCD15, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD557, 16'hB411, 16'hAB8E, 16'hFE9B, 16'hFEDC, 16'hCCD3, 16'h7985, 16'hAB8F, 16'hD556, 16'hCD15, 16'hCD15, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC4D4, 16'hC493, 16'hCCD4, 16'hC4D4, 16'hC4D4, 16'hC494, 16'hC494, 16'hC494, 16'hC4D4, 16'hC4D4, 16'hC493, 16'hC493, 16'hB410, 16'hC452, 16'hCC93, 16'hABD0, 16'hB3D0, 16'hABCF, 16'hC4D4, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515,
        16'hC4D4, 16'hC4D4, 16'h7A89, 16'h938D, 16'hD555, 16'hA3CF, 16'h7248, 16'h9B8F, 16'hB452, 16'h934E, 16'hB492, 16'h9BCF, 16'hC4D4, 16'h7249, 16'hABCF, 16'hCCD3, 16'hC492, 16'h6207, 16'hAC93, 16'hBD15, 16'hBD15, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'hBD14, 16'hBD15, 16'hB4D4, 16'hB514, 16'hBD15, 16'hBD15, 16'hC556, 16'h834D, 16'hAC92, 16'hD5D7, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hDDD8, 16'hE619, 16'hFEDC, 16'hF69B, 16'hEE19, 16'hCD15, 16'hE5D8, 16'hCD14, 16'hEE5A, 16'hBC52, 16'hF6DC, 16'hFF1E, 16'hFEDD, 16'hF69B, 16'hDD98, 16'hDD97, 16'hDD97, 16'hD557, 16'hD556, 16'hAC11, 16'hC4D4, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hC494, 16'hCCD5, 16'hCCD5, 16'hCD15, 16'hCCD5, 16'hD516, 16'hA38F, 16'hABCF, 16'hDD97, 16'h8A8A, 16'hC492, 16'h8B0C, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hD556, 16'hCCD4, 16'hC493, 16'hD516, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516,
        16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'hBC52, 16'hA34D, 16'hFE9B, 16'hFEDC, 16'hE5D8, 16'h8A49, 16'h92CA, 16'hCD14, 16'hD556, 16'hCD15, 16'hD516, 16'hD516, 16'hD516, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hCCD4, 16'hC493, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC494, 16'hC494, 16'hC494, 16'hC4D4, 16'hC4D4, 16'hC493, 16'hC494, 16'hB411, 16'hB411, 16'hCC93, 16'hB411, 16'hB3CF, 16'hABD0, 16'hBC93, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D4, 16'hCD15, 16'h8B0C, 16'h72CA, 16'hCD14, 16'h9B8E, 16'h7248, 16'h938E, 16'hBCD3, 16'h938E, 16'hB493, 16'h8B4D, 16'hC4D4, 16'h8B4D, 16'h8ACB, 16'hCCD3, 16'hCCD3, 16'h934C, 16'h834D, 16'hBD15, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'hB514, 16'hBD15, 16'hB4D5, 16'hB4D4, 16'hBD15, 16'hBD15, 16'hC556, 16'h9C10, 16'h8B8D, 16'hDE18, 16'hDE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hF69B, 16'hD515, 16'hABCF, 16'hDDD8, 16'hE5D8, 16'hCD15, 16'hE619, 16'hB452, 16'hFF1D, 16'hFF1D, 16'hFEDD,
        16'hE619, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD15, 16'hABD0, 16'hCCD5, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hCD15, 16'hCD15, 16'hC4D4, 16'hC494, 16'hCCD5, 16'hCCD5, 16'hCD15, 16'hCCD5, 16'hD515, 16'h92CC, 16'hC4D4, 16'hDD56, 16'h8249, 16'hC493, 16'h82CB, 16'hCD15, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hD556, 16'hCD15, 16'hBC52, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'hCCD4, 16'h9B0B, 16'hF69B, 16'hF6DC, 16'hFE9B, 16'hABCF, 16'h81C6, 16'hBC11, 16'hDD56, 16'hCCD5, 16'hD516, 16'hD516, 16'hD516, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hCCD5, 16'hC494, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC494, 16'hC494, 16'hC4D4, 16'hC4D4, 16'hC493, 16'hC494, 16'hBC52, 16'hABD0, 16'hCC93, 16'hBC52, 16'hAB8F,
        16'hB3D0, 16'hBC93, 16'hCD15, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D4, 16'hCD15, 16'hAC10, 16'h61C6, 16'hC513, 16'h9B8E, 16'h7249, 16'h938E, 16'hC514, 16'h938E, 16'hB492, 16'h8B4D, 16'hBC93, 16'hB451, 16'h69C7, 16'hBC51, 16'hCCD3, 16'hBC51, 16'h7248, 16'hAC93, 16'hBD15, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'hBD14, 16'hBD15, 16'hBCD5, 16'hB4D4, 16'hBD15, 16'hBD15, 16'hBD56, 16'hAC93, 16'h7289, 16'hD5D7, 16'hD5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF6DC, 16'hC492, 16'hBC93, 16'hEEDB, 16'hFF1D, 16'hDDD7, 16'hDDD8, 16'hDD97, 16'hCD15, 16'hFF5E, 16'hFEDD, 16'hFEDC, 16'hDD98, 16'hCD15, 16'hCD16, 16'hCD15, 16'hCD56, 16'hC493, 16'hABD0, 16'hCD15, 16'hC4D5, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC4D4, 16'hC4D4, 16'hCCD5, 16'hCCD5, 16'hCCD5, 16'hCD15, 16'hC4D4, 16'h7A49, 16'hEDD8, 16'hD556, 16'h92CB, 16'hCCD3, 16'h82CB, 16'hCCD5, 16'hD516, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hCD15, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD16, 16'hCD15, 16'hBC52,
        16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'hD516, 16'hD516, 16'hD516, 16'hD515, 16'h928A, 16'hEE59, 16'hFEDC, 16'hFEDC, 16'hDD96, 16'h8186, 16'h9B0D, 16'hDD56, 16'hCD15, 16'hCD15, 16'hD516, 16'hD516, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hCCD5, 16'hCCD4, 16'hC494, 16'hCCD4, 16'hC4D4, 16'hC494, 16'hC494, 16'hC494, 16'hC4D4, 16'hC4D4, 16'hC493, 16'hC493, 16'hC493, 16'hA38F, 16'hC452, 16'hC493, 16'hA34E, 16'hB411, 16'hB452, 16'hCD15, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D4, 16'hC515, 16'hB452, 16'h6A07, 16'hBCD3, 16'h9B8E, 16'h7249, 16'h7ACB, 16'hC514, 16'hAC10, 16'hB452, 16'h938E, 16'hA411, 16'hCD15, 16'h82CB, 16'h930C, 16'hCCD3, 16'hCCD4, 16'h934C, 16'h8B8E, 16'hBD15, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD5, 16'hBCD5, 16'hB4D4,
        16'hBD15, 16'hBD15, 16'hBD16, 16'hB514, 16'h6A08, 16'hC596, 16'hD5D7, 16'hF79D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF1D,
        16'hBC93, 16'hCD56, 16'hFF9F, 16'hF71D, 16'hF71C, 16'hD597, 16'hE619, 16'hC4D4, 16'hE619, 16'hFF5E, 16'hFEDD, 16'hF69B, 16'hD556, 16'hCD15, 16'hCD15, 16'hC515, 16'hCD15, 16'hB452, 16'hB452, 16'hCD15, 16'hC4D5, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hC4D4, 16'hC4D4, 16'hCCD5, 16'hCCD5, 16'hCCD5, 16'hD516, 16'hABD0, 16'h9B4D, 16'hFE9B, 16'hDD96, 16'h8ACA, 16'hCD14, 16'h7249, 16'hC4D4, 16'hD516, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC4D4, 16'hCD15, 16'hCD16, 16'hCD15, 16'hCCD5, 16'hD516, 16'hCD16, 16'hCD15, 16'hCD16, 16'hD516, 16'hBC52, 16'hCD15, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'hD556, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'h928A, 16'hDDD7, 16'hFF1D, 16'hF69B, 16'hF69B, 16'hAB8E, 16'h79C7, 16'hC493, 16'hD516, 16'hC4D4, 16'hD516, 16'hD516, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hCCD5, 16'hCCD4, 16'hCCD4, 16'hC493, 16'hCCD4, 16'hC4D4,
        16'hC494, 16'hC493, 16'hC493, 16'hC4D4, 16'hC4D4, 16'hC493, 16'hC493, 16'hC493, 16'hB3D0, 16'hB3D0, 16'hCCD3, 16'h9B4E, 16'hBC11, 16'hB452, 16'hC515, 16'hC4D5, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D4, 16'hC515, 16'hC4D4, 16'h6A07, 16'hAC10, 16'h9B8E, 16'h7249, 16'h8B4C, 16'hC515, 16'hAC11, 16'hAC51, 16'h9BD0, 16'h9BCF, 16'hCD55, 16'hAC51, 16'h6A08, 16'hBC51, 16'hCCD3, 16'hB451, 16'h6A49, 16'hB493, 16'hBCD4, 16'hB4D4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'hB4D4, 16'hBD15, 16'hB4D4, 16'hB4D4, 16'hBD15, 16'hBD15, 16'hBD15, 16'h7A8B, 16'hB4D3, 16'hE618, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hCD55, 16'hDE19, 16'hFFDF, 16'hFFDF, 16'hEE9B, 16'hFF9E, 16'hCD56, 16'hEE5A, 16'hB3D0, 16'hF69B, 16'hFF1D, 16'hFEDD, 16'hF65B, 16'hCD15, 16'hCD15, 16'hC4D4, 16'hC4D4, 16'hCD15, 16'hABD0, 16'hBC93, 16'hCD15, 16'hC4D4, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hCCD5, 16'hCCD4, 16'hCCD4, 16'hC4D4, 16'hC4D4, 16'hCCD5, 16'hCCD5, 16'hCCD5, 16'hD515, 16'h8ACC, 16'hAC10, 16'hFEDC, 16'hDD97, 16'h92CB, 16'hD514, 16'h6186, 16'hB452, 16'hD556, 16'hCD15, 16'hCD15,
        16'hCD15, 16'hC4D4, 16'hCD15, 16'hCD16, 16'hCD15, 16'hCCD5, 16'hD516, 16'hCD16, 16'hCD15, 16'hCD16, 16'hD516, 16'hBC52, 16'hCCD4, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD16, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hDD57, 16'h9ACC, 16'hD596, 16'hFF5E, 16'hF69C, 16'hFEDC, 16'hDD56, 16'h7944, 16'hA38E, 16'hDD56, 16'hC4D4, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hCCD5, 16'hCCD4, 16'hCCD4, 16'hC493, 16'hC493, 16'hC4D4, 16'hC494, 16'hC493, 16'hC493, 16'hC4D4, 16'hC4D4, 16'hC4D3, 16'hC493, 16'hC493, 16'hBC52, 16'hA34E, 16'hCCD3, 16'h9B4D, 16'hB410, 16'hB451, 16'hCD15, 16'hC4D4, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC514, 16'hC514, 16'hC514, 16'hCD15, 16'h7A8A, 16'h9B8E, 16'hAC10, 16'h61C7, 16'h9BCF, 16'hC515, 16'hBC93, 16'h9BCF, 16'hAC51, 16'h9BCF, 16'hC514, 16'hC4D4, 16'h7249, 16'hA38E, 16'hCCD3, 16'hCCD3, 16'h82CB,
        16'h9BD0, 16'hBD14, 16'hB4D4, 16'hBCD4, 16'hB4D4, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'hBCD4, 16'hB4D4, 16'hBD14, 16'hB4D4, 16'hB4D4, 16'hBD15, 16'hBD15, 16'hBD16, 16'h938E, 16'h93CF, 16'hDE19, 16'hDE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hE69B, 16'hFF9E, 16'hCD15, 16'hE619, 16'hBC52, 16'hFF1D, 16'hFF1D, 16'hFEDC, 16'hE619, 16'hC4D5, 16'hCD15, 16'hBCD4, 16'hC515, 16'hC515, 16'hA38F, 16'hC4D4, 16'hC515, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hC4D4, 16'hCCD5, 16'hCCD4, 16'hC4D4, 16'hC4D4, 16'hCCD4, 16'hCCD5, 16'hCCD5, 16'hCD15, 16'hCD15, 16'h8249, 16'hD515, 16'hFEDC, 16'hDD97, 16'h8289, 16'hD514, 16'h7208, 16'hABD0, 16'hD556, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC4D4, 16'hCD15, 16'hCD16, 16'hCD15, 16'hCCD5, 16'hCD15, 16'hCD16, 16'hCD16, 16'hCD16, 16'hD556, 16'hC493, 16'hC4D4, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hDD97, 16'hA34E, 16'hC514, 16'hFFDF, 16'hFF1D, 16'hF69B, 16'hF65A, 16'hAB8E, 16'h7186, 16'hCD14, 16'hCD15, 16'hCD15,
        16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hCCD5, 16'hCCD4, 16'hCCD4, 16'hC4D4, 16'hC493, 16'hC4D4, 16'hC493, 16'hC493, 16'hC493, 16'hC493, 16'hC4D4, 16'hC4D4, 16'hC493, 16'hC493, 16'hC493, 16'h9B4E, 16'hBC52, 16'hA34E, 16'hABD0, 16'hB411, 16'hCD15, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC514, 16'hC514, 16'hC514, 16'hCD15, 16'h8B4D, 16'h7ACA, 16'hA3CF, 16'h5103, 16'h9BCF, 16'hC514, 16'hBCD3, 16'h938E, 16'hB492, 16'h8B4D, 16'hC514, 16'hC514, 16'h9BCF, 16'h7A49, 16'hC492, 16'hCCD4, 16'hB451, 16'h6A89, 16'hB4D3, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'hB4D4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'hBD14, 16'hBCD4, 16'hB4D4, 16'hBD15, 16'hBD15, 16'hBD16, 16'hA411, 16'h7B0C, 16'hD5D8, 16'hDDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hF75D, 16'hEF1C, 16'hC4D4, 16'hD556, 16'hCD15, 16'hFF1E, 16'hFEDD, 16'hFEDC, 16'hDDD8, 16'hC4D4, 16'hCD15, 16'hC4D4, 16'hCD15, 16'hBCD3, 16'hA390, 16'hC4D5, 16'hC4D4, 16'hC4D5, 16'hC4D5, 16'hC4D5, 16'hCCD5, 16'hCCD5, 16'hCCD5, 16'hCCD4, 16'hC4D4, 16'hCCD5, 16'hCCD5, 16'hCCD5, 16'hCD15,
        16'hC4D4, 16'h8ACB, 16'hEE19, 16'hFE9C, 16'hDD97, 16'h8249, 16'hD515, 16'h7A49, 16'h9B8E, 16'hD516, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hCD15, 16'hCD16, 16'hCD15, 16'hCCD5, 16'hCD15, 16'hCD16, 16'hCD16, 16'hCD16, 16'hD556, 16'hC4D4, 16'hC493, 16'hD516, 16'hCD16, 16'hCD16, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'hD556, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD557, 16'hDD98, 16'hB411, 16'hBC51, 16'hFFDF, 16'hFF9F, 16'hFF1D, 16'hFEDC, 16'hEE18, 16'h8249, 16'hA38E, 16'hD556, 16'hC4D4, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hCCD5, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hC493, 16'hC494, 16'hC493, 16'hC493, 16'hC493, 16'hC493, 16'hC4D4, 16'hC4D4, 16'hC493, 16'hC493, 16'hC493, 16'hAB8F, 16'hABCF, 16'h9B4E, 16'hABCF, 16'hB411, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D4, 16'hCD15, 16'h9BCF, 16'h82CA, 16'hA3CE, 16'h50C2, 16'h9B8E,
        16'hC514, 16'hC514, 16'h938E, 16'hB452, 16'h8B4D, 16'hBCD3, 16'hC514, 16'hBCD3, 16'h6A08, 16'hABCF, 16'hCCD3, 16'hCCD4, 16'h7ACA, 16'h9BD0, 16'hBD14, 16'hB4D4, 16'hBCD4, 16'hB493, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'hB4D4, 16'hBCD4, 16'hB4D4, 16'hBD15, 16'hBD15, 16'hBD16, 16'hAC93, 16'h830C, 16'hC596, 16'hD5D6, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'hFFDF, 16'hDE59, 16'hCD15, 16'hBC93, 16'hDDD8, 16'hFF1E, 16'hFEDC, 16'hF69B, 16'hD597, 16'hC4D5, 16'hCD15, 16'hBC93, 16'hCD15, 16'hBC92, 16'hAC11, 16'hC4D5, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hCCD5, 16'hCCD5, 16'hCCD4, 16'hC4D4, 16'hCCD5, 16'hCCD5, 16'hCCD5, 16'hCD15, 16'hB411, 16'h930D, 16'hF65A, 16'hFE9B, 16'hDD97, 16'h7A48, 16'hD555, 16'h828A, 16'h82CB, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD16, 16'hCD15, 16'hCCD5, 16'hCD15, 16'hCD15, 16'hC4D4, 16'hCD15, 16'hCD16, 16'hCD16, 16'hCD16, 16'hD516, 16'hCCD5, 16'hBC93, 16'hCD16, 16'hCD16, 16'hCD16, 16'hD516, 16'hD516, 16'hD556, 16'hD556, 16'hD556, 16'hD516, 16'hD516, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hDD97, 16'hD557, 16'hD556,
        16'hD515, 16'hB3CF, 16'h9B4D, 16'hFF9E, 16'hF75D, 16'hD555, 16'hCD14, 16'hC4D3, 16'h930C, 16'h5904, 16'hCCD4, 16'hCD15, 16'hCD15, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hCCD5, 16'hCCD5, 16'hCCD4, 16'hCCD4, 16'hC493, 16'hC493, 16'hC493, 16'hC493, 16'hC493, 16'hC493, 16'hC4D4, 16'hC4D4, 16'hC493, 16'hC493, 16'hC493, 16'hBC52, 16'hA38E, 16'hAB8F, 16'hABD0, 16'hB410, 16'hC4D4, 16'hC515, 16'hC515, 16'hCD15, 16'hCD15, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D4, 16'hCD15, 16'hB451, 16'h7289, 16'hABCE, 16'h5102, 16'h9BCE, 16'hC514, 16'hC514, 16'h9BCF, 16'hAC51, 16'h938E, 16'hAC52, 16'hC514, 16'hC514, 16'h938E, 16'h7A8A, 16'hCCD3, 16'hD4D3, 16'hABCF, 16'h7ACB, 16'hBCD4, 16'hB4D4, 16'hBCD4, 16'hB4D3, 16'hB4D4, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'hB4D4, 16'hBCD4, 16'hB4D4, 16'hB515, 16'hBD15, 16'hBD16, 16'hAC93, 16'h830D, 16'hB514, 16'hDDD8, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1D, 16'hDE18, 16'hFFDF, 16'hCD96, 16'hD597, 16'hBC92, 16'hE619, 16'hFF1D, 16'hFEDC, 16'hEE5A, 16'hCD55, 16'hC4D4, 16'hC515, 16'hBC93, 16'hCD15, 16'hB411, 16'hAC11, 16'hCD15, 16'hC4D4,
        16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hCCD4, 16'hC4D4, 16'hC4D4, 16'hCCD4, 16'hCCD4, 16'hCCD5, 16'hD515, 16'h930D, 16'hBC92, 16'hFE9B, 16'hFE9B, 16'hE5D8, 16'h8289, 16'hDD56, 16'h930C, 16'h828A, 16'hC4D4, 16'hD556, 16'hCD15, 16'hCD56, 16'hCD15, 16'hCCD5, 16'hCD16, 16'hCD16, 16'hCCD5, 16'hCD15, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hD515, 16'hC493, 16'hCD16, 16'hCD16, 16'hCD16, 16'hD516, 16'hD516, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD557, 16'hD556, 16'hBC52, 16'hABCF, 16'hA34E, 16'h8A8A, 16'h9A8A, 16'h8249, 16'hD596, 16'hDDD7, 16'hD4D3, 16'hBC10, 16'h9B0C, 16'h8ACA, 16'h59C6, 16'h934D, 16'hC493, 16'hC493, 16'hCD15, 16'hD515, 16'hD516, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCCD5, 16'hCCD4, 16'hC4D3, 16'hC493, 16'hC493, 16'hC493, 16'hC493, 16'hC493, 16'hC493, 16'hC4D4, 16'hC493, 16'hC493, 16'hC493, 16'hC493, 16'hA38E, 16'h9B0C, 16'hABCF, 16'hBC51, 16'hC4D4, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15,
        16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D4, 16'hCD15, 16'hBCD3, 16'h6A48, 16'hA3CE, 16'h6185, 16'h938E, 16'hC514, 16'hC514, 16'hAC10, 16'hA410, 16'hA410, 16'h9C10, 16'hC514, 16'hBD14, 16'hB492, 16'h61C7, 16'hB451, 16'hCCD3, 16'hC492, 16'h7A8A, 16'hAC51, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'hB4D3, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB514, 16'hB4D4, 16'hB514, 16'hBD15, 16'hBD16, 16'hB4D4, 16'h8B4D, 16'hA451, 16'hDDD8, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'hEEDB, 16'hFFDF, 16'hC514, 16'hD596, 16'hBC52, 16'hF6DC, 16'hFF1D, 16'hF69B, 16'hE619, 16'hCD56, 16'hC515, 16'hC515, 16'hBC93, 16'hCD15, 16'hABD0, 16'hBC53, 16'hC515, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hCCD4, 16'hC4D4, 16'hC4D4, 16'hCCD4, 16'hCCD4, 16'hCCD5, 16'hCD15, 16'h8A8B, 16'hD556, 16'hFE9B, 16'hFEDC, 16'hEE5A, 16'h92CB, 16'hE596, 16'h930C, 16'h934D, 16'hBC92, 16'hD556, 16'hCD15, 16'hCD56, 16'hCD15, 16'hCCD5, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hD516, 16'hC493, 16'hCD15, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'hD556, 16'hD556,
        16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCCD4, 16'h9B0C, 16'h5000, 16'h6144, 16'h7A49, 16'h828A, 16'h7A08, 16'h79C7, 16'hCD14, 16'hD556, 16'hC4D3, 16'hAB8E, 16'hA34D, 16'h6986, 16'h4840, 16'h4104, 16'h6A07, 16'h7248, 16'h9B4D, 16'hB411, 16'hBC92, 16'hCCD4, 16'hD556, 16'hCD15, 16'hCD15, 16'hC4D5, 16'hCCD4, 16'hC4D4, 16'hC493, 16'hC493, 16'hC493, 16'hC493, 16'hC493, 16'hC493, 16'hC4D4, 16'hC4D3, 16'hC493, 16'hC493, 16'hC493, 16'hABCF, 16'h8ACA, 16'hABCF, 16'hBC51, 16'hC4D4, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC514, 16'h7ACA, 16'h934C, 16'h6185, 16'h93CE, 16'hC514, 16'hC4D4, 16'hB492, 16'h9B8E, 16'hA410, 16'h93CE, 16'hC514, 16'hBCD3, 16'hC514, 16'h830C, 16'h934D, 16'hCCD3, 16'hC492, 16'h934C, 16'h8B4D, 16'hBD14, 16'hB4D4, 16'hB4D4, 16'hB493, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'hB4D4, 16'hB514, 16'hB4D4, 16'hB4D4, 16'hBD15, 16'hBD15, 16'hB4D4, 16'h93CF, 16'h93CF, 16'hDDD8,
        16'hD5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hF79E, 16'hFFDF, 16'hC514, 16'hD597, 16'hBC92, 16'hFF1D,
        16'hFEDC, 16'hEE9B, 16'hE619, 16'hCD15, 16'hC515, 16'hC4D4, 16'hBC93, 16'hCD15, 16'hA3D0, 16'hBC94, 16'hC4D5, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hCCD4, 16'hC4D4, 16'hC4D4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCD15, 16'hC4D4, 16'h828A, 16'hEE19, 16'hFE9B, 16'hFF1D, 16'hF71C, 16'h8ACA, 16'hDD96, 16'hA38E, 16'h9B8E, 16'hA3CF, 16'hD556, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD16, 16'hCD15, 16'hCD15, 16'hD516, 16'hCD16, 16'hCD16, 16'hD516, 16'hD556, 16'hC4D4, 16'hCCD4, 16'hD556, 16'hD516, 16'hD516, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD516, 16'hD516, 16'hD557, 16'hC494, 16'h92CB, 16'h930D, 16'hABD0, 16'hBC52, 16'hC494, 16'hD516, 16'hCCD4, 16'h9249, 16'hEE9A, 16'hFFDF, 16'hFF9E, 16'hF71C, 16'hEE59, 16'hDD97, 16'hCD14, 16'h7A89, 16'h5185, 16'h5185, 16'h48C0, 16'h69C7, 16'h7208, 16'h8ACB, 16'hAC10, 16'hC493, 16'hD515, 16'hCD15, 16'hCCD4, 16'hC4D4, 16'hC493, 16'hC493, 16'hC493, 16'hC493, 16'hC493, 16'hC493, 16'hC4D3, 16'hC4D3, 16'hC493,
        16'hC493, 16'hC493, 16'hBC51, 16'h8248, 16'hA38F, 16'hBC52, 16'hC4D3, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D4, 16'hCD15, 16'h9B8E, 16'h82CA, 16'h5985, 16'h9BCE, 16'hC514, 16'hBCD4, 16'hBCD3, 16'h938E, 16'hAC51, 16'h938E, 16'hC514, 16'hBCD4, 16'hBD14, 16'hA451, 16'h6A07, 16'hBC91, 16'hC492, 16'h934C, 16'h7A8A, 16'hB493, 16'hBCD4, 16'hB4D4, 16'hB493, 16'hB4D4, 16'hBCD4, 16'hB4D4, 16'hB4D4, 16'hB514, 16'hB4D4, 16'hB4D4, 16'hB515, 16'hBD56, 16'hBD15, 16'h93CF, 16'h834E, 16'hCD96, 16'hD596, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hDE18, 16'hFFDF, 16'hFF9E, 16'hC4D4, 16'hCD14, 16'hCD15, 16'hFF1D, 16'hF6DC, 16'hEE5A, 16'hE5D8, 16'hCD15, 16'hC515, 16'hC4D4, 16'hBC93, 16'hC4D4, 16'hA3D0, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hCCD4, 16'hC4D4, 16'hC4D4, 16'hCCD4, 16'hCCD5, 16'hCCD4, 16'hCD15, 16'hB411, 16'hA38E, 16'hFE9B, 16'hFEDC, 16'hFF5E, 16'hFF5E, 16'h9B4C, 16'hE618, 16'hB452, 16'hA3CE, 16'h934D, 16'hD556, 16'hD516, 16'hD516, 16'hD556, 16'hCD15, 16'hCD15, 16'hCD56, 16'hCD15, 16'hCD15, 16'hD516,
        16'hCD16, 16'hCD16, 16'hD516, 16'hD556, 16'hCCD5, 16'hC4D4, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD516, 16'hCCD5, 16'hDD57, 16'hD516, 16'hD515, 16'hDD56, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hE597, 16'h9249, 16'hD5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hFF1D, 16'hFEDC, 16'hE5D7, 16'h8208, 16'hBC51, 16'hC452, 16'h9B8E, 16'h7A8A, 16'h6A07, 16'h5102, 16'h6A07, 16'hA3CF, 16'hCCD4, 16'hD515, 16'hCCD4, 16'hC494, 16'hC493, 16'hC493, 16'hC493, 16'hC493, 16'hC493, 16'hC4D3, 16'hC4D3, 16'hC4D4, 16'hC493, 16'hC493, 16'hC453, 16'h8249, 16'hA34E, 16'hC493, 16'hC493, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D4, 16'hCD15, 16'hA3D0, 16'h6A07, 16'h61C6, 16'h8B4C, 16'hC514, 16'hBCD3, 16'hBCD4, 16'h938E, 16'hA410, 16'h938D, 16'hBD14, 16'hBCD4, 16'hBCD4, 16'hBCD3, 16'h6A49, 16'hA3CE, 16'hABCF, 16'h7A8A, 16'hAC10, 16'hB493, 16'hBCD4, 16'hBCD4, 16'hB493, 16'hB493,
        16'hBCD4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hACD4, 16'hC556, 16'h93D0, 16'h838E, 16'hC515, 16'hD596, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'hE659, 16'hFFDF, 16'hEF1C, 16'hBC93, 16'hC4D4, 16'hD596, 16'hFF1D, 16'hF69C, 16'hEE5A, 16'hDDD7, 16'hC515, 16'hC515, 16'hC4D5, 16'hC4D4, 16'hBC93, 16'hA3D0, 16'hC515, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D5, 16'hC4D4, 16'hC4D4, 16'hCCD5, 16'hC4D4, 16'hC4D4, 16'hD515, 16'h9B4E, 16'hB411, 16'hFE9B, 16'hF69B, 16'hFF9E, 16'hFFDF, 16'h9B4D, 16'hDDD7, 16'hB493, 16'hBC92, 16'h934D, 16'hC4D4, 16'hD556, 16'hD516, 16'hD556, 16'hCD15, 16'hCD15, 16'hCD16, 16'hCD16, 16'hCD15, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'hD516, 16'hCCD4, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD557, 16'hDD56, 16'hC452, 16'hDD56, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hE597, 16'hA30D, 16'hC514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hFEDD, 16'hFEDD, 16'hFEDC, 16'hABCF, 16'h930C, 16'hE597, 16'hDD56, 16'hD515, 16'hCCD4, 16'hBC51, 16'h8ACC, 16'h71C7,
        16'h7A08, 16'hB410, 16'hCCD4, 16'hC4D4, 16'hC494, 16'hC494, 16'hC494, 16'hC494, 16'hC493, 16'hC4D3, 16'hC4D4, 16'hC4D4, 16'hC494, 16'hC493, 16'hCCD4, 16'h828A, 16'h8ACC, 16'hC493, 16'hC493, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D4, 16'hCD15, 16'hAC11, 16'h5985, 16'h6A07, 16'h8B0C, 16'hC4D4, 16'hBCD3, 16'hC514, 16'h9BCF, 16'hA410, 16'h8B4D, 16'hB4D3, 16'hBD14, 16'hBCD4, 16'hC514, 16'h8B8D, 16'h8B0B, 16'h7A89, 16'h830C, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'hBCD4, 16'hB493, 16'hAC51, 16'hBCD4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'h9411, 16'hBD56, 16'h9C52, 16'h8BCF, 16'hB4D3, 16'hDDD7, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hEEDB, 16'hFFDF, 16'hEEDB, 16'hBC52, 16'hB411, 16'hEE19, 16'hFEDD, 16'hF69B, 16'hE619, 16'hD597, 16'hC515, 16'hC515, 16'hC4D4, 16'hC4D4, 16'hAC12, 16'hAC11, 16'hC515, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D5, 16'hC4D4, 16'hC4D4, 16'hC4D5, 16'hCD15, 16'hCD15, 16'hCD15, 16'h82CC, 16'hA38E, 16'hA38E, 16'hCCD3, 16'hDE18, 16'hE65A, 16'h938E, 16'h930B, 16'hA38E,
        16'hCD14, 16'h9B8D, 16'hAC11, 16'hDD57, 16'hD516, 16'hD556, 16'hD516, 16'hCD15, 16'hCD16, 16'hCD16, 16'hCD15, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD556, 16'hD556, 16'hCCD4, 16'hD516, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hDD57, 16'hDD57, 16'hDD57, 16'hBC10, 16'hD4D5, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hE598, 16'hBBD0, 16'hABCF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5D, 16'hFF1C, 16'hFF1D, 16'hEE19, 16'h79C7, 16'hBC11, 16'hE557, 16'hD516, 16'hD516, 16'hDD56, 16'hD515, 16'hCCD4, 16'hBC11, 16'h9B0D, 16'hABCF, 16'hC493, 16'hBC52, 16'hCCD4, 16'hC494, 16'hC494, 16'hC494, 16'hC4D4, 16'hC4D4, 16'hCCD4, 16'hCCD4, 16'hC494, 16'hCCD4, 16'hA34E, 16'h92CB, 16'hC493, 16'hC493, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC515, 16'hC515, 16'hC515, 16'hC4D4, 16'hC515, 16'hB452, 16'h5985, 16'h6207, 16'h830C, 16'hC4D4, 16'hBCD3, 16'hBD14, 16'hA410, 16'h9BCF, 16'h938D, 16'hAC92, 16'hBD14,
        16'hBCD4, 16'hBD14, 16'hA450, 16'h59C5, 16'h7289, 16'hAC92, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBC93, 16'h9BCF, 16'hBCD4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB514, 16'hB4D4, 16'hB515, 16'hA452, 16'hB515, 16'hACD3, 16'h8BD0, 16'hAC92, 16'hDDD7, 16'hDE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE659, 16'hF75D, 16'hFFDF, 16'hEF1C, 16'hB410, 16'hA3CF, 16'hF69B, 16'hFEDC, 16'hF69B, 16'hE619, 16'hD556, 16'hC4D4, 16'hCD15, 16'hC4D4, 16'hC4D4, 16'hA3D1, 16'hB452, 16'hC4D5, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hCCD5, 16'hC4D4, 16'hCCD4, 16'hCD15, 16'hC4D3, 16'hA38F, 16'h828A, 16'h6186, 16'h8249, 16'h79C7, 16'h928A, 16'hA30C, 16'hBC93, 16'hA3D0, 16'hB451, 16'hC514, 16'hBC92, 16'hBC51, 16'h934D, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD15, 16'hCD16, 16'hD556, 16'hCD15, 16'hD515, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD15, 16'hD515, 16'hD557, 16'hD556, 16'hD556, 16'hD556, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hE597, 16'hBC11, 16'hB3D0, 16'hE598, 16'hDD57, 16'hDD97, 16'hDD57, 16'hDD57, 16'hDD97, 16'hDD97, 16'hE598, 16'hCC93, 16'h9ACB, 16'hFF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFF9E, 16'hFF1D, 16'hFEDC, 16'hFF1D, 16'hCCD4, 16'h6903, 16'hDD15, 16'hDD56, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD515, 16'hCCD4, 16'hD4D5, 16'hA38E, 16'hC452, 16'hCCD4, 16'hC494, 16'hC4D4, 16'hC4D4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hC493, 16'hCCD4, 16'hB3D0, 16'h828A, 16'hC493, 16'hC493, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC515, 16'hC4D5, 16'hC515, 16'hBC93, 16'h61C7, 16'h61C5, 16'h82CB, 16'hBCD3, 16'hBC93, 16'hBCD4, 16'hAC51, 16'h9B8E, 16'h9B8E, 16'hA410, 16'hC514, 16'hBCD4, 16'hBCD4, 16'hAC92, 16'h5185, 16'h8B4E, 16'hBCD4, 16'hB4D3, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'h8B4E, 16'hAC52, 16'hBCD5, 16'hB4D4, 16'hB514, 16'hBD14, 16'hACD4, 16'hB515, 16'hA493, 16'hA493, 16'hBD55, 16'h9410, 16'h9C11, 16'hD5D7, 16'hD5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hEF5E, 16'hEF5D, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDDD8, 16'hFF9E, 16'hFFDF, 16'hE69B, 16'hB3D0, 16'hBC93, 16'hFEDC, 16'hF69C, 16'hEE5A, 16'hE5D9, 16'hD556, 16'hC4D4, 16'hC515, 16'hC4D4, 16'hC4D4, 16'hAC11, 16'hBC93, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hCD14, 16'hA3D0,
        16'h8ACC, 16'h5944, 16'h50C3, 16'h5104, 16'h938E, 16'hB451, 16'hD596, 16'hEEDB, 16'hFF9F, 16'hD597, 16'hC514, 16'hE659, 16'hABCF, 16'hCD14, 16'h9B4D, 16'hC4D4, 16'hDD57, 16'hD556, 16'hD556, 16'hCD15, 16'hCD16, 16'hD556, 16'hCD15, 16'hCCD4, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD515, 16'hD556, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hE597, 16'hCC93, 16'h9249, 16'hE557, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD98, 16'hDD97, 16'hDD97, 16'hE598, 16'hDD16, 16'h89C7, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hFEDC, 16'hFEDD, 16'hFEDB, 16'h930C, 16'h9B4D, 16'hE597, 16'hDD56, 16'hD516, 16'hD516, 16'hD516, 16'hD516, 16'hD515, 16'hD515, 16'hD515, 16'hBC11, 16'hAB8F, 16'hCCD5, 16'hC4D4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hC494, 16'hCCD4, 16'hBC11, 16'h8249, 16'hC493, 16'hC493, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC515, 16'hC515,
        16'hC4D4, 16'h6A08, 16'h5143, 16'h8B4C, 16'hBCD3, 16'hBC93, 16'hBCD3, 16'hB492, 16'h938D, 16'h9BCF, 16'h9BCF, 16'hC514, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'h830C, 16'h938F, 16'hBCD4, 16'hB4D3, 16'hB4D4, 16'hB4D4, 16'hBCD4, 16'hBCD4, 16'h938F, 16'h9BD0, 16'hBD15, 16'hB4D4, 16'hB514, 16'hB515, 16'hB4D4, 16'hB515, 16'hACD4, 16'h9C51, 16'hBD56, 16'h8B8F, 16'hA452, 16'hD5D7, 16'hCD55, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DC, 16'hD65A,
        16'hCDD9, 16'hCDD9, 16'hCE1A, 16'hDE5B, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hDE19, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'h81C7, 16'hCD15, 16'hFF1D, 16'hF69C, 16'hEE5A, 16'hE5D8, 16'hD556, 16'hC4D4, 16'hC515, 16'hC4D5, 16'hC4D4, 16'hB411, 16'hBC93, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hCD14, 16'hB411, 16'h82CC, 16'h48C2, 16'h4882, 16'h7ACB, 16'h8ACC, 16'hAC10, 16'hFEDC, 16'hFF1D, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hAC10, 16'hEEDC, 16'hC4D3, 16'hDDD7, 16'hABCF, 16'hA38F, 16'hDD97, 16'hD556, 16'hD556, 16'hD556, 16'hCD16, 16'hD556, 16'hD556, 16'hB3D1, 16'hD516, 16'hD556, 16'hD556, 16'hD557, 16'hD557, 16'hDD56, 16'hD515, 16'hD556, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hE557, 16'hDD16, 16'h91C7, 16'hCC93, 16'hE598,
        16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'h9A0A, 16'hD618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF1D, 16'hFEDC, 16'hFF1D, 16'hEE19, 16'h7A07, 16'hB411, 16'hE597, 16'hDD56, 16'hDD56, 16'hDD56, 16'hDD16, 16'hD556, 16'hD515, 16'hD515, 16'hCCD4, 16'h8A8A, 16'hC493, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hC493, 16'h7A08, 16'hBC52, 16'hC494, 16'hCD15, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC515, 16'hCD14, 16'h82CB, 16'h48C1, 16'hB451, 16'hBCD4, 16'hBC93, 16'hBC93, 16'hBCD3, 16'h938E, 16'hAC10, 16'h938E, 16'hBD14, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hB493, 16'hAC52, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hB493, 16'hB4D4, 16'hBCD4, 16'h9C10, 16'h830D, 16'hBCD4, 16'hB4D4, 16'hB4D4, 16'hB515, 16'hB4D4, 16'hB515, 16'hB515, 16'h9410, 16'hBD55, 16'h9410, 16'h9C51, 16'hDE18, 16'hCD14, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1D, 16'hCDDA, 16'hC5D9, 16'hCDDA, 16'hCE1A, 16'hCDD9, 16'hC5D9, 16'hCE1A, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'hE65A, 16'hFFDF, 16'hFFDF, 16'hDE18, 16'h9249, 16'hE5D8, 16'hFF1D, 16'hF69B, 16'hEE19, 16'hE5D8, 16'hCD15, 16'hC4D4, 16'hC515, 16'hC4D5, 16'hC4D4, 16'hAC11,
        16'hBC94, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hCD15, 16'hAC11, 16'h6187, 16'h3800, 16'h6A08, 16'hAC10, 16'hD555, 16'hA34E, 16'hD555, 16'hFF1D, 16'hF71C, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h9B8D, 16'hE618, 16'hBC92, 16'hD555, 16'hC492, 16'hA34E, 16'hD556, 16'hD557, 16'hD556, 16'hD556, 16'hCD16, 16'hD556, 16'hDD97, 16'hA34E, 16'hC493, 16'hDD97, 16'hD556, 16'hDD57, 16'hDD57, 16'hDD57, 16'hD556, 16'hD556, 16'hDD57, 16'hDD57, 16'hDD97, 16'hDD97, 16'hDD97, 16'hE597, 16'hE597, 16'hE597, 16'hE557, 16'hB34D, 16'hB34E, 16'hE597, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hED98, 16'hA2CC, 16'hCD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF1D, 16'hFEDC, 16'hFF1D, 16'hD555, 16'h5000, 16'hD514, 16'hDD57, 16'hDD56, 16'hDD56, 16'hDD56, 16'hDD56, 16'hDD56, 16'hD515, 16'hD515, 16'h9B0C, 16'hABCF, 16'hD515, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'h8A8A, 16'hC452, 16'hCCD4, 16'hCD15,
        16'hCD16, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC515, 16'hCD15, 16'h8B0C, 16'h4000, 16'hA410, 16'hBCD4, 16'hB493, 16'hB493, 16'hBCD4, 16'h9B8E, 16'hA410, 16'h9B8E, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hAC92, 16'hB493, 16'hBCD4, 16'hAC52, 16'h82CC, 16'hAC92, 16'hBD15, 16'hB4D4, 16'hB515, 16'hB4D4, 16'hB4D5, 16'hBD55, 16'h9411, 16'hB515, 16'h9C52, 16'h93D0, 16'hE69A, 16'hC4D3, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79F, 16'hCDDA, 16'hCE1A, 16'hCE1A, 16'hC5DA, 16'hCDDA, 16'hCE1A, 16'hCE1A, 16'hC5D9, 16'hD65B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9B, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hBD14, 16'h928A, 16'hEE9A, 16'hFF1D, 16'hF69B, 16'hE619, 16'hDDD8, 16'hCD56, 16'hC4D4, 16'hC515, 16'hC515, 16'hC4D4, 16'hA38F, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hCD15, 16'hA3D0, 16'h4000, 16'h5986, 16'h9B8E, 16'hCCD4, 16'hD556, 16'hCCD4, 16'h8A08, 16'hE619, 16'hFF1D, 16'hFF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB451, 16'hDD96, 16'hBC92, 16'hDE18, 16'hCD14, 16'hABCF, 16'hC492, 16'hDD97, 16'hD556, 16'hDD57, 16'hD556, 16'hD556, 16'hDD97, 16'hBC11, 16'hA34E, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD57, 16'hD556,
        16'hDD97, 16'hDD97, 16'hDD97, 16'hDD97, 16'hE598, 16'hE597, 16'hE598, 16'hE597, 16'hED98, 16'hCC52, 16'hB34D, 16'hD493, 16'hEDD9, 16'hE598, 16'hEDD9, 16'hE598, 16'hE598, 16'hE598, 16'hEDD9, 16'hC411, 16'hBC51, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFF1D, 16'hFF1D, 16'hFF1C, 16'hBC92, 16'h8248, 16'hDD56, 16'hE557, 16'hDD56, 16'hDD56, 16'hDD56, 16'hDD56, 16'hD516, 16'hDD56, 16'hC452, 16'h8208, 16'hCCD3, 16'hCCD5, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'h92CB, 16'hBC51, 16'hCCD4, 16'hCD15, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC515, 16'hC515, 16'hCD15, 16'h9B4E, 16'h50C1, 16'h9B8E, 16'hBCD4, 16'hB493, 16'hB493, 16'hBCD4, 16'h9BCF, 16'hA3CF, 16'h938E, 16'hB493, 16'hBCD4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hB493, 16'hB493, 16'hBCD4, 16'hB493, 16'h830D, 16'h9BD0, 16'hBD15, 16'hB4D4, 16'hB514, 16'hB4D4, 16'hB4D4, 16'hBD16,
        16'h9C11, 16'hACD4, 16'hACD3, 16'h838E, 16'hEF1C, 16'hC4D3, 16'hD5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hCDD9, 16'hCE1A, 16'hCE1A, 16'hC5DA, 16'hCDDA, 16'hCDD9, 16'hCDDA, 16'hCDD9, 16'hCE1A, 16'hF79F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65A, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hB4D3,
        16'h7987, 16'hF69B, 16'hFF1D, 16'hF65B, 16'hE5D8, 16'hDDD8, 16'hCD15, 16'hC4D5, 16'hC515, 16'hC515, 16'hC4D4, 16'hAC11, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hCD15, 16'hA38F, 16'h3800, 16'h830C, 16'hBC92, 16'hD555, 16'hD556, 16'hD556, 16'hB411, 16'hAB8E, 16'hFF1C, 16'hFF1C, 16'hFF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC555, 16'hD555, 16'hDDD7, 16'hD555, 16'hD514, 16'hC492, 16'hA38E, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD57, 16'hD556, 16'hDD97, 16'hCCD4, 16'h8A09, 16'hD516, 16'hDD98, 16'hDD57, 16'hDD57, 16'hDD97, 16'hE597, 16'hDD57, 16'hDD57, 16'hE597, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hED98, 16'hD493, 16'hC3D0, 16'hCC11, 16'hE557, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hE598, 16'hEDD9, 16'hD4D5, 16'hAB0C, 16'hFF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFF1D, 16'hFF1D, 16'hFEDC, 16'hA3CE, 16'h8A8A, 16'hDD55, 16'hDD57, 16'hDD56, 16'hDD57, 16'hDD56, 16'hDD56, 16'hDD56, 16'hDD56, 16'h8A8B, 16'h9B4E,
        16'hD515, 16'hCCD5, 16'hCD15, 16'hCCD5, 16'hCCD5, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'h92CB, 16'hB410, 16'hCCD4, 16'hCD15, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC515, 16'hCD15, 16'hA3CF, 16'h6185, 16'h8B0C, 16'hB493, 16'hBC93, 16'hBC93, 16'hBCD4, 16'hA411, 16'h9B8E, 16'h9B8E, 16'hAC92, 16'hBD14, 16'hB4D4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'hBCD4, 16'hB4D3, 16'hAC52, 16'hBCD4, 16'hBCD4, 16'h934E, 16'h834D, 16'hB4D4, 16'hB515, 16'hB514, 16'hB4D4, 16'hB4D4, 16'hBD16, 16'hA452, 16'hA492, 16'hBD55, 16'h7B0C, 16'hEEDC, 16'hDE18, 16'hC4D3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1D, 16'hC5D9, 16'hCE1A, 16'hCE1A, 16'hCDDA, 16'hCDDA, 16'hCDDA, 16'hCDDA, 16'hCDDA, 16'hCDD9, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hAC51, 16'h9B0D, 16'hF6DC, 16'hFF1D, 16'hEE5A, 16'hE5D8, 16'hDD98, 16'hC515, 16'hC4D5, 16'hC515, 16'hC4D5, 16'hC4D4, 16'hB452, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hCCD4, 16'h8ACC, 16'h7A8A, 16'h6A07, 16'hB451, 16'hCCD4, 16'hCD15, 16'hD515, 16'hD556, 16'hB3D0, 16'hB451, 16'hFF1D, 16'hF71C, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hAC51, 16'hDDD7, 16'hB491, 16'hDE17, 16'hD514, 16'hBC92, 16'hC493, 16'hE598, 16'hDD97,
        16'hDD97, 16'hD556, 16'hDD97, 16'hDD56, 16'h924A, 16'hBBD1, 16'hE598, 16'hE557, 16'hE597, 16'hE598, 16'hE598, 16'hE597, 16'hDD57, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hED98, 16'hE557, 16'hCC11, 16'hDD15, 16'hC3CF, 16'hF5D9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hE557, 16'hAA4A, 16'hE659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFF1D, 16'hFF1D, 16'hFE9B, 16'h9B4D, 16'h928A, 16'hE596, 16'hE597, 16'hDD57, 16'hDD57, 16'hDD57, 16'hDD56, 16'hDD57, 16'hBC11, 16'h7186, 16'hCCD4, 16'hD515, 16'hCD15, 16'hD515, 16'hCD15, 16'hCD15, 16'hCCD4, 16'hCCD4, 16'hA30D, 16'hB3D0, 16'hCCD4, 16'hCD15, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC515, 16'hCD15, 16'hABD0, 16'h6186, 16'h7A89, 16'hAC51, 16'hBCD4, 16'hBCD3, 16'hBCD4, 16'hAC52, 16'h9B8E, 16'h9B8E, 16'hA410, 16'hBD14, 16'hB4D4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4,
        16'hB4D4, 16'hA411, 16'hB4D3, 16'hBCD4, 16'hA410, 16'h7ACC, 16'hA451, 16'hBD15, 16'hB514, 16'hB515, 16'hB4D4, 16'hBD15, 16'hACD3, 16'h9411, 16'hBD55, 16'h730C, 16'hDE9B, 16'hEF1C, 16'hB451, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hCDDA, 16'hCE1A, 16'hCE1A, 16'hCDDA, 16'hCDDA, 16'hCDDA, 16'hCDDA, 16'hCDDA, 16'hCE1A, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE18, 16'hF71D, 16'hFFDF, 16'hFF9F, 16'hA3D0, 16'hB410, 16'hFF5E, 16'hFF1D, 16'hEE5A, 16'hE5D8, 16'hDDD8, 16'hC515, 16'hC4D5, 16'hC4D4, 16'hC515, 16'hBC93, 16'hA38F, 16'hC4D4, 16'hC4D4, 16'hC4D5, 16'hC4D4, 16'h8ACC, 16'hA3CF, 16'hBC93, 16'h7249, 16'hC4D3, 16'hCCD4, 16'hD555, 16'hD515, 16'hDD56, 16'h9B0C, 16'hC4D3, 16'hFF5D, 16'hFF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAC51, 16'hD555, 16'hBC92, 16'hEE9A, 16'hC4D2, 16'hD513, 16'hAB8F, 16'hE598, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD57, 16'hE597, 16'hB38F, 16'hA2CB, 16'hD4D5, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hE598, 16'hED98, 16'hED98, 16'hED98, 16'hE598, 16'hEDD9, 16'hD411, 16'hE597, 16'hD4D3, 16'hD452, 16'hF61A, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hF5D9, 16'hC38F, 16'hD595, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5E,
        16'hFF1E, 16'hFE9B, 16'hA34D, 16'h92CB, 16'hE597, 16'hE598, 16'hDD57, 16'hE557, 16'hDD57, 16'hDD57, 16'hDD56, 16'h8248, 16'hABCF, 16'hDD56, 16'hCD15, 16'hD515, 16'hD515, 16'hD515, 16'hCD15, 16'hD4D4, 16'hA34D, 16'hBC11, 16'hD515, 16'hCD15, 16'hCD16, 16'hCD16, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC515, 16'hCD15, 16'hB451, 16'h69C6, 16'h7A48, 16'hA3D0, 16'hBCD4, 16'hBC93, 16'hBCD3, 16'hB493, 16'h9B8E, 16'hA3CF, 16'h9BCF, 16'hBD14, 16'hB4D4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'hBCD4, 16'hA411, 16'hAC92, 16'hBD15, 16'hAC51, 16'h830D, 16'h93D0, 16'hBD15, 16'hB514, 16'hB515, 16'hB4D4, 16'hB515, 16'hB4D4, 16'h9411, 16'hB555, 16'h7B0C, 16'hD659, 16'hFF9F, 16'hB410, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF69C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hD61B, 16'hCDD9, 16'hCE1A, 16'hCE1A, 16'hCE1A, 16'hCDDA, 16'hCDDA, 16'hC5D9, 16'hD69B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD5D7, 16'hF75D, 16'hFFDF, 16'hFF9E, 16'hB411, 16'hABCF, 16'hFF1D, 16'hFF1D, 16'hEE1A, 16'hE5D8, 16'hDD97, 16'hC515, 16'hC4D5, 16'hC4D4, 16'hC515, 16'hBC93, 16'hABD0, 16'hC4D5, 16'hC4D4, 16'hCD15, 16'hAC11, 16'hA3D0, 16'hD515, 16'hAC11, 16'h5986, 16'hC4D3, 16'hCCD4, 16'hD555, 16'hD555, 16'hD555, 16'h92CC, 16'hE619, 16'hFF5D, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'hB450, 16'hD514, 16'hE659, 16'hD5D7, 16'hDDD7, 16'hB492, 16'hD4D4, 16'hE5D8, 16'hE598, 16'hE598, 16'hDD57, 16'hE598, 16'hCC52, 16'hC38F, 16'hB38F, 16'hED98, 16'hE598, 16'hE598, 16'hED98, 16'hED98, 16'hED98, 16'hE597, 16'hEDD8, 16'hED98, 16'hED99, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hE556, 16'hCC52, 16'hF6DC, 16'hB34D, 16'hE515, 16'hF61A, 16'hEDD9, 16'hF5D9, 16'hEDD9, 16'hF5D9, 16'hDCD5, 16'hC3CF, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hF69B, 16'h9B0C, 16'h9249, 16'hDD15, 16'hE598, 16'hE597, 16'hE597, 16'hDD57, 16'hE597, 16'hBC11, 16'h6000, 16'hCC93, 16'hD556, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD4D4, 16'hA30D, 16'hABD0, 16'hD4D5, 16'hCD15, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hBC52, 16'h69C7, 16'h934D, 16'h934D, 16'hBCD3, 16'hBCD3, 16'hBCD3,
        16'hBCD3, 16'h938D, 16'hA3CF, 16'h938E, 16'hBCD4, 16'hB4D4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hAC52, 16'hA452, 16'hBD15, 16'hAC92, 16'h8B4E, 16'h938F, 16'hBD14, 16'hBD14, 16'hB515, 16'hB4D4, 16'hB515, 16'hB515, 16'h9411, 16'hB515, 16'h7B4D, 16'hC596, 16'hFFDF, 16'hBCD4, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hCE1A, 16'hC5D9, 16'hCE1A, 16'hCE1A, 16'hCDDA, 16'hC5D9, 16'hC5D9, 16'hEF5D, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD596, 16'hF75D, 16'hFFDF, 16'hEF1C, 16'h9B4D, 16'hB411, 16'hFF5E, 16'hFF1D, 16'hEE19, 16'hE5D8, 16'hDD97, 16'hC515, 16'hC4D4, 16'hC4D4, 16'hC515, 16'hBC93, 16'hABD0, 16'hC4D5, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC515, 16'hCD15, 16'h934E, 16'h6A08, 16'hC4D3, 16'hCD14, 16'hD556, 16'hD556, 16'hCD15, 16'h8A8A, 16'hEE5A, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDE, 16'hB451, 16'hC492, 16'hD5D7, 16'hFF5D, 16'hC513, 16'hE659, 16'hAB4D, 16'hE598, 16'hE5D8, 16'hE5D8, 16'hE598, 16'hE598, 16'hD4D5, 16'hCBD0, 16'hCC10, 16'hCC52, 16'hF5D9, 16'hEDD8, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hDD15, 16'hE516, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hF5D9, 16'hC30E, 16'hE5D8, 16'hFF1D, 16'hB30E, 16'hE516, 16'hFE5A, 16'hEDD9, 16'hEDD9, 16'hF5D9,
        16'hF5D9, 16'hBB0E, 16'hEE5A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF1C, 16'hB411, 16'h8144, 16'hC452, 16'hE598, 16'hE598, 16'hDD97, 16'hE597, 16'hE556, 16'h8A49, 16'h8ACB, 16'hDD56, 16'hD556, 16'hD556, 16'hD516, 16'hD515, 16'hD4D4, 16'hA30C, 16'hB410, 16'hD515, 16'hD516, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hBC93, 16'h69C6, 16'hA410, 16'h82CB, 16'hAC51, 16'hBCD4, 16'hB493, 16'hBCD4, 16'h9B8E, 16'hA3CF, 16'h938D, 16'hB4D3, 16'hBCD4, 16'hB4D4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hB493, 16'h9BD0, 16'hBD15, 16'hB4D3, 16'h93CF, 16'h8B4E, 16'hB4D4, 16'hBD15, 16'hBD15, 16'hB4D5, 16'hB515, 16'hBD15, 16'h9C52, 16'hA493, 16'h838E, 16'hB4D4, 16'hFFDF, 16'hD618, 16'hCD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71D, 16'hD61A, 16'hCDD9, 16'hC5D9, 16'hC5D9, 16'hCE1A, 16'hEF1D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD5D7, 16'hFF9E, 16'hFFDF, 16'hEEDB, 16'hAB4E, 16'hC492, 16'hFF5E, 16'hFEDC, 16'hE619, 16'hE5D8, 16'hDD97, 16'hC4D5, 16'hC4D4, 16'hC4D4, 16'hC515, 16'hBC52, 16'hA3CF, 16'hC515, 16'hC4D4, 16'hC4D4, 16'hC4D5, 16'hC4D5, 16'hC4D4, 16'h8ACC, 16'h7A8A,
        16'hCCD4, 16'hCD15, 16'hD556, 16'hDD56, 16'hC493, 16'h930C, 16'hF6DC, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9B, 16'h92CA, 16'hB450, 16'hFFDF, 16'hD596, 16'hDDD7, 16'hCD14, 16'hB38F, 16'hF619, 16'hEDD9, 16'hEDD9, 16'hE5D8, 16'hEDD8, 16'hCC11, 16'hDC94, 16'hBB4E, 16'hE556, 16'hF5D9, 16'hEDD9, 16'hEDD9, 16'hF5D9, 16'hED98, 16'hD452, 16'hED98, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hF61A, 16'hDCD4, 16'hCC51, 16'hFFDF, 16'hEEDB, 16'hB2CC, 16'hE516, 16'hFE1A, 16'hF61A, 16'hF5D9, 16'hF61A, 16'hD453, 16'hC451, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hD556, 16'h7900, 16'hB38F, 16'hE557, 16'hEDD8, 16'hEDD8, 16'hE598, 16'hD4D4, 16'h6000, 16'hBC52, 16'hDD97, 16'hD556, 16'hD556, 16'hD556, 16'hD4D4, 16'h9ACB, 16'hB410, 16'hD515, 16'hD556, 16'hCD56, 16'hD556, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD15,
        16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC4D4, 16'h71C7, 16'hAC10, 16'h934D, 16'h9B8E, 16'hC4D4, 16'hBCD3, 16'hBCD4, 16'hAC10, 16'h9BCE, 16'h938E, 16'hB493, 16'hBCD4, 16'hB4D4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'h9BD0, 16'hB4D4, 16'hBCD4, 16'h9C10, 16'h938F, 16'hA452, 16'hBD15, 16'hB515, 16'hB515, 16'hB515, 16'hBD55, 16'hA452, 16'h9C93, 16'h8C10, 16'hA451, 16'hFFDF, 16'hEEDC, 16'hC514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hEF1D, 16'hE6DC, 16'hEF1D, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD96, 16'hFF9E, 16'hFFDF, 16'hDE59, 16'hB3CF, 16'hC492, 16'hFF5E, 16'hF6DC, 16'hE5D8, 16'hE5D8, 16'hD597, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'hC515, 16'hBC52, 16'hA38F, 16'hCD15, 16'hC4D4, 16'hC4D5, 16'hC4D5, 16'hCD15, 16'hBC52, 16'h92CB, 16'h8ACC, 16'hC493, 16'hD555, 16'hD556, 16'hDD97, 16'hBC11, 16'hC492, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD96, 16'hA34C, 16'hF71C, 16'hFFDF, 16'hBC10, 16'hE5D8, 16'hBC52, 16'hD493, 16'hF61A, 16'hEDD9, 16'hEDD9, 16'hF619, 16'hDCD5, 16'hCC12, 16'hE515, 16'hBB4D, 16'hF5D8, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF61A, 16'hE516, 16'hD453, 16'hF61A, 16'hF5DA, 16'hF5D9, 16'hF5D9,
        16'hF5DA, 16'hF5D9, 16'hF5DA, 16'hF5D9, 16'hC30E, 16'hE598, 16'hFFDF, 16'hF71C, 16'hD493, 16'hCB90, 16'hED57, 16'hFE1A, 16'hFE1A, 16'hF599, 16'hC34F, 16'hF6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hB411, 16'h9249, 16'hB3CF, 16'hD515, 16'hE598, 16'hF619, 16'hBC11, 16'h8249, 16'hD555, 16'hDD56, 16'hD556, 16'hD556, 16'hDD15, 16'hA34D, 16'hB3D0, 16'hD515, 16'hCD16, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCCD4, 16'h7208, 16'hA410, 16'hB451, 16'h7A8A, 16'hBCD3, 16'hBCD4, 16'hBCD4, 16'hB451, 16'h9B8D, 16'h9B8E, 16'hAC52, 16'hBCD4, 16'hB4D4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBD14, 16'h9C11, 16'hAC92, 16'hBD15, 16'h9C11, 16'h8B8E, 16'h93CF, 16'hBD15, 16'hB515, 16'hB4D4, 16'hB515, 16'hB515, 16'hA493, 16'h9C93, 16'h9C52, 16'h93CF, 16'hF75D, 16'hFF9F, 16'hBCD3,
        16'hF79D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hCD96, 16'hFF9E, 16'hFFDF, 16'hDDD8, 16'hC493, 16'hC493, 16'hFF5E, 16'hF6DC, 16'hE5D9, 16'hE5D8, 16'hDD97, 16'hC4D4, 16'hC4D5,
        16'hC4D4, 16'hC515, 16'hBC52, 16'hA38F, 16'hCD15, 16'hC4D4, 16'hC515, 16'hC4D5, 16'hD515, 16'hABCF, 16'h9B4D, 16'h9B0C, 16'hC4D3, 16'hD556, 16'hD556, 16'hDD97, 16'hAB8F, 16'hD515, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC4D3, 16'hB410, 16'hFFDF, 16'hF71C, 16'hC492, 16'hEE19, 16'hB34E, 16'hDD15, 16'hF61A, 16'hF5D9, 16'hEDD9, 16'hF5D9, 16'hCC10, 16'hE5D8, 16'hDCD4, 16'hCB8E, 16'hF5D9, 16'hF61A, 16'hF5DA, 16'hF61A, 16'hFE1A, 16'hDC94, 16'hD453, 16'hF61A, 16'hF61A, 16'hF5DA, 16'hF61A, 16'hF61A, 16'hF5D9, 16'hF61A, 16'hED57, 16'hC34F, 16'hF6DB, 16'hFFDF, 16'hFF9E, 16'hDD97, 16'hBB4F, 16'hDC52, 16'hED97, 16'hF5D9, 16'hE4D5, 16'hD451, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hF75D, 16'hF75D, 16'hFF5E, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hEE5A, 16'hBC92, 16'hA2CB, 16'h9A8A, 16'hC451, 16'hDCD4, 16'h7103, 16'hA34D, 16'hDD56, 16'hDD56, 16'hDD56, 16'hDD56,
        16'h9B0C, 16'hB410, 16'hD515, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD56, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'h8289, 16'hA3CF, 16'hCD14, 16'h828A, 16'hBC92, 16'hC514, 16'hBCD4, 16'hB493, 16'h934D, 16'h9BCE, 16'hA411, 16'hBCD4, 16'hB4D4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBD14, 16'hAC52, 16'hA411, 16'hBD15, 16'hA451, 16'h93CF, 16'h938F, 16'hB514, 16'hB515, 16'hB4D4, 16'hB515, 16'hB555, 16'hACD3, 16'h9C52, 16'hA493, 16'h8B4D, 16'hE6DB, 16'hFFDF, 16'hCD55, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hCD96, 16'hFF9E, 16'hFFDF, 16'hD596, 16'hC4D3, 16'hCD15, 16'hFF5E, 16'hF69B, 16'hE5D9, 16'hE5D9, 16'hD597, 16'hC4D4, 16'hC4D5, 16'hC4D4, 16'hC515, 16'hB452, 16'hA38F, 16'hCD15, 16'hC4D4, 16'hC515, 16'hC515, 16'hD515, 16'h930D, 16'hB410, 16'h9B0D, 16'hCCD3, 16'hDD56, 16'hDD56, 16'hDD56, 16'hAB4D, 16'hEE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hC4D3, 16'hE658, 16'hFFDF, 16'hEE5A, 16'hC411, 16'hDD55, 16'hBB8F, 16'hE516, 16'hFE1A, 16'hF5D9, 16'hF5D9, 16'hED56, 16'hCC11,
        16'hFE9C, 16'hCC93, 16'hC38F, 16'hF5D8, 16'hF65B, 16'hF61A, 16'hF619, 16'hFE19, 16'hDCD4, 16'hD452, 16'hE557, 16'hFE5B, 16'hF61A, 16'hF61A, 16'hF5D9, 16'hF5D9, 16'hF61A, 16'hE516, 16'hC38F, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFF5D, 16'hD4D5, 16'hC30D, 16'hCB4F, 16'hD3D1, 16'hD3D0, 16'hEDD8, 16'hEE9A, 16'hD555, 16'hC411, 16'hB34E, 16'h928A, 16'h92CB, 16'h92CB, 16'h9B0C, 16'hBC92, 16'hCD15, 16'hDE18, 16'hF6DC, 16'hFF5D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF71C, 16'hE659, 16'hC514, 16'hC492, 16'hC451, 16'h81C7, 16'hBC11, 16'hDD56, 16'hD556, 16'hDD56, 16'hA30D, 16'hB3D0, 16'hD515, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'h930C, 16'h934D, 16'hD555, 16'h8B0C, 16'hAC51, 16'hCD15, 16'hC514, 16'hBCD4, 16'h934C, 16'h9B8E, 16'h9BCF, 16'hBCD4, 16'hB4D4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hB493, 16'h9BD0, 16'hBD15, 16'hAC52, 16'h93CF, 16'h8B4E,
        16'hAC93, 16'hB515, 16'hB4D5, 16'hB515, 16'hB515, 16'hB515, 16'h9C51, 16'hA4D3, 16'h938F, 16'hD618, 16'hFFDF, 16'hD618, 16'hCDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD55,
        16'hFF9E, 16'hFF9F, 16'hC514, 16'hC4D3, 16'hC4D4, 16'hFF5E, 16'hF69B, 16'hE5D9, 16'hE5D9, 16'hDD97, 16'hC4D4, 16'hC4D5, 16'hC4D4, 16'hC515, 16'hB452, 16'hA34E, 16'hCD15, 16'hCCD5, 16'hCCD5, 16'hCD15, 16'hC4D4, 16'h71C7, 16'hD514, 16'h9B4D, 16'hBC52, 16'hDD56, 16'hDD96, 16'hD515, 16'hAB8E, 16'hF75C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE18, 16'hEEDB, 16'hFFDF, 16'hF71C, 16'hD514, 16'hDCD4, 16'hC34E, 16'hE4D4, 16'hF5D8, 16'hF5D9, 16'hFE19, 16'hE4D5, 16'hCC52, 16'hFEDD, 16'hDD15, 16'hBB0C, 16'hE515, 16'hF61A, 16'hFE5A, 16'hFE5B, 16'hFE5B, 16'hED98, 16'hCC11, 16'hDC94, 16'hF5D9, 16'hFE5B, 16'hFE5A, 16'hF61A, 16'hF61A, 16'hFE5B, 16'hE556, 16'hCC93, 16'hF6DC, 16'hFF5E, 16'hFF5E, 16'hF69B, 16'hE5D8, 16'hEE19, 16'hEDD8, 16'hE4D4, 16'hCBCF, 16'hB209, 16'hA1C6, 16'hB34D, 16'hB3CF, 16'hB38E, 16'hB38E, 16'h9ACB, 16'hAB8E, 16'hA34C, 16'hA34C, 16'hAB8D, 16'hAB8D, 16'hB3CF, 16'hC4D3, 16'hEE5A,
        16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hDD97, 16'h89C7, 16'hCCD3, 16'hDD56, 16'hDD56, 16'hAB8E, 16'hB3D0, 16'hCCD4, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'h934D, 16'h7ACA, 16'hD596, 16'h9B8E, 16'h82CB, 16'hB452, 16'hCD55, 16'hC514, 16'h9B8E, 16'h9B8E, 16'h9BCF, 16'hBCD4, 16'hB4D4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'h9C10, 16'hB4D4, 16'hAC93, 16'h93CF, 16'h938F, 16'h9C11, 16'hBD15, 16'hB514, 16'hB515, 16'hB515, 16'hBD56, 16'h9411, 16'h8C10, 16'hA492, 16'hCD96, 16'hFFDF, 16'hE6DB, 16'hBD14, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD96, 16'hF75D, 16'hFF5E, 16'hC514, 16'hD5D7, 16'hC514, 16'hFF5E, 16'hEE5A, 16'hE619, 16'hE619, 16'hDD97, 16'hC4D4, 16'hC4D5, 16'hC4D4, 16'hC515, 16'hBC52, 16'h9B4E, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hB451, 16'h828B, 16'hEE18, 16'h9B0C, 16'hBC52, 16'hE597, 16'hE597, 16'hD515, 16'hC452, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hEEDB, 16'hEE9A, 16'hFFDF, 16'hFFDF, 16'hF6DC, 16'hEE18, 16'hD451, 16'hCB8F, 16'hE4D4, 16'hF598, 16'hFE19, 16'hE4D5, 16'hD4D4, 16'hFF1D, 16'hEE1A, 16'hD411, 16'hCB8E, 16'hD452, 16'hE4D4, 16'hED98, 16'hF5D9, 16'hED56, 16'hDC94, 16'hD453, 16'hD452, 16'hDC93, 16'hEDD8, 16'hF619, 16'hE555, 16'hED98, 16'hEE9B, 16'hE5D9, 16'hE597, 16'hF6DB, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hEE19, 16'hCC52, 16'hDD55, 16'hE619, 16'hF71C, 16'hF6DB, 16'hDD56, 16'hCC51, 16'hC410, 16'hA34C, 16'h930B, 16'h8B0B, 16'h7A89, 16'h8B0B, 16'hA34C, 16'hA30C, 16'h9B0B, 16'h9ACB, 16'hBC51, 16'hDDD7, 16'hEEDC, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC514, 16'h81C6, 16'hCCD4, 16'hE597, 16'hB38F, 16'hBC10, 16'hD515, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD15, 16'hA3CF, 16'h7248, 16'hD596, 16'hB451, 16'hA38E, 16'h82CC, 16'hA3D0, 16'hCD55, 16'h9BCF, 16'h9B8E, 16'h938E, 16'hB4D4, 16'hBCD4, 16'hBCD4,
        16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'hBCD4, 16'h9C10, 16'hAC93, 16'hB4D4, 16'h93D0, 16'hA411, 16'h93D0, 16'hBD15, 16'hB514, 16'hB515, 16'hB515, 16'hBD56, 16'h9411, 16'h7B8E, 16'hB514, 16'hC555, 16'hFFDF, 16'hF79E, 16'hBCD3, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD5D7, 16'hFF5E, 16'hF71D, 16'hCD15, 16'hD5D7, 16'hCD15, 16'hFF5E, 16'hEE5A, 16'hE619, 16'hE619, 16'hDD97, 16'hC4D4, 16'hC4D5, 16'hC4D5, 16'hC515, 16'hBC93, 16'h9B8E, 16'hCD15, 16'hCD15, 16'hCD15, 16'hD516, 16'hABD0, 16'h9B4E, 16'hFE9B, 16'hAB8E, 16'hC492, 16'hE5D8, 16'hE5D8, 16'hCCD4, 16'hDDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5D, 16'hE597, 16'hCC10, 16'hCB4E, 16'hDC11, 16'hECD5, 16'hD3D0, 16'hD452, 16'hEDD9, 16'hF65A, 16'hEE19, 16'hE5D8, 16'hD4D3, 16'hD4D3, 16'hE555, 16'hF69A, 16'hFF9F, 16'hF71D, 16'hE5D8, 16'hCCD3, 16'hD4D4, 16'hE597, 16'hE5D8, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE59, 16'hDD97, 16'hF75D, 16'hFFDF, 16'hF71D, 16'hDE18, 16'hABCF,
        16'h8A89, 16'h71C6, 16'h5102, 16'h5944, 16'h4902, 16'h4944, 16'h4903, 16'h4943, 16'h5185, 16'h61C6, 16'h7208, 16'h7A89, 16'h930A, 16'h8A48, 16'hAB8D, 16'hCD14, 16'hF6DC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hB450, 16'h7986, 16'hDD15, 16'hB3CF, 16'hB3CF, 16'hD515, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD16, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD56, 16'hB451, 16'h7206, 16'hD556, 16'hB492, 16'h934D, 16'hBC93, 16'h6186, 16'hBCD3, 16'hB452, 16'h934D, 16'h938E, 16'hB4D3, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'hB4D4, 16'hBD14, 16'hA452, 16'hAC52, 16'hBD15, 16'h93CF, 16'h9C10, 16'h8B4E, 16'hB514, 16'hB515, 16'hB515, 16'hB515, 16'hBD96, 16'h9C92, 16'h838E, 16'hBD96, 16'hC556, 16'hF75D, 16'hFFDF, 16'hBD14, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD5D8, 16'hFF5E, 16'hEEDB, 16'hCD55, 16'hC514, 16'hCD55, 16'hFF5E, 16'hEE5A, 16'hE619, 16'hE619, 16'hDD97, 16'hC4D5, 16'hC515, 16'hC515, 16'hCD15, 16'hBC93, 16'h9B4E, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'h8A8A, 16'hBC93, 16'hFEDC, 16'hB410, 16'hCCD3, 16'hE5D8, 16'hE5D8, 16'hD515, 16'hF6DC, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hEEDB, 16'hDDD8, 16'hCD55, 16'hBCD3, 16'hBCD3, 16'hC514, 16'hDDD7, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5D, 16'hEE5A, 16'hEDD8, 16'hDD96, 16'hEE5A, 16'hEE9A, 16'hEE99, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFFDF, 16'hFF5E, 16'hCD55, 16'h8A08, 16'h6800, 16'h4800, 16'h5104, 16'h5985, 16'h4944, 16'h4103, 16'h4904, 16'h4103, 16'h5184, 16'h5985, 16'h5184, 16'h4944, 16'h4103, 16'h4944, 16'h4944, 16'h6A07, 16'h7208, 16'h7A06, 16'hABCE, 16'hE5D8, 16'hFF5E, 16'hFF9F, 16'hFFDF, 16'hFF5E, 16'hB410, 16'h9ACB, 16'hA30C, 16'hBC10, 16'hD4D4, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD16, 16'hCD56, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD56, 16'hBC92, 16'h69C5,
        16'hCD14, 16'hCD14, 16'h8289, 16'hC514, 16'h8B4D, 16'h8B4D, 16'hB492, 16'h8B4C, 16'h938D, 16'hB4D3, 16'hBD14, 16'hBCD4, 16'hB4D4, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hBD14, 16'hAC93, 16'hA411, 16'hBD15, 16'h9C10, 16'hA411, 16'h8B8E, 16'hACD4, 16'hB515, 16'hB515, 16'hB515, 16'hC597, 16'hA493, 16'h734D, 16'hBD96, 16'hCD97, 16'hE69A, 16'hFFDF, 16'hCDD7, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD5D7, 16'hF71D, 16'hE65A, 16'hCD15, 16'hCD55, 16'hCD15, 16'hFF5E, 16'hEE1A, 16'hE619, 16'hE619, 16'hDD97, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC493, 16'h930D, 16'hCCD5, 16'hCD15, 16'hCD16, 16'hC4D4, 16'h79C7, 16'hE5D8, 16'hFF1D, 16'hC493, 16'hC452, 16'hF619, 16'hEDD8, 16'hE5D7, 16'hEE59, 16'hFF1D, 16'hEE19, 16'hB411, 16'h9ACB, 16'hA2CB, 16'h9249, 16'hA2CC, 16'hAB0C, 16'h9A8A, 16'h8986, 16'h9A89, 16'hABCF, 16'hDDD7, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5D, 16'hEEDB, 16'hF6DB, 16'hEE18, 16'hA30C, 16'h6800, 16'h6985, 16'h69C6, 16'h61C6, 16'h5944, 16'h4880, 16'h48C2, 16'h5144, 16'h4944, 16'h4944, 16'h4944, 16'h5184, 16'h4944, 16'h4944, 16'h5144, 16'h4944, 16'h4944, 16'h4103, 16'h38C2, 16'h5185, 16'h7207, 16'h9ACA, 16'hD4D3, 16'hFF1C, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hBC92, 16'h6800, 16'hB3CF, 16'hD4D4, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD16, 16'hD556, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD16, 16'hC492, 16'h71C6, 16'hC514, 16'hD555, 16'h8289, 16'hC4D3, 16'hC514, 16'h6A49, 16'hA3CF, 16'h938E, 16'h8B4D, 16'hAC92, 16'hBD14, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'hB4D4, 16'hB514, 16'hB4D4, 16'h93D0, 16'hB4D4, 16'hA452, 16'hA451, 16'h8B8E, 16'hA452, 16'hBD56, 16'hAD15, 16'hB515, 16'hBD97, 16'hAD14, 16'h7B8E, 16'hBD96, 16'hD619, 16'hD5D7, 16'hFFDF, 16'hE69A, 16'hCDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hEE9B, 16'hE659, 16'hC514, 16'hD5D7, 16'hCD55, 16'hFF1D, 16'hEE5A, 16'hE619, 16'hE619, 16'hD597, 16'hC4D5, 16'hC515, 16'hC4D4, 16'hC4D4, 16'hC4D4, 16'h930D, 16'hCCD4, 16'hCD15, 16'hD556, 16'hB411,
        16'h930C, 16'hF65A, 16'hFF1D, 16'hDD97, 16'hC452, 16'hD515, 16'hC452, 16'hBC10, 16'hE5D7, 16'hE597, 16'hB38E, 16'hA30C, 16'hAB4D, 16'hA34D, 16'hAB4D, 16'hC451, 16'hCC51, 16'hCC51, 16'hDD14, 16'hDD55, 16'hD555, 16'hC452, 16'hCCD4, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hDD97, 16'hD4D4, 16'hEE19, 16'hCC92, 16'h8944, 16'h7144, 16'h7A07, 16'h7186, 16'h71C6, 16'h58C0, 16'h69C6, 16'h8B0B, 16'h8B0B, 16'h82CA, 16'h7289, 16'h6A48, 16'h6207, 16'h59C6, 16'h5144, 16'h4944, 16'h4944, 16'h5144, 16'h5985, 16'h5185, 16'h4103, 16'h38C2, 16'h4103, 16'h5184, 16'h8A89, 16'hDD14, 16'hEE9A, 16'hFF9F, 16'hFFDF, 16'hFF5D, 16'hA38E, 16'hAB4D, 16'hD4D4, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556,
        16'hD556, 16'hD556, 16'hCD16, 16'hD556, 16'hD556, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD16, 16'hC4D3, 16'h7A07, 16'hC4D3, 16'hD556, 16'h7A49, 16'hBC92, 16'hD596, 16'h938E, 16'h7A8A, 16'h9BCF, 16'h834C, 16'hAC92, 16'hBD14, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hBCD4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'h9BD0, 16'hACD3, 16'hAC92, 16'h9C10, 16'hA451, 16'h93D0, 16'hBD55, 16'hB515, 16'hACD4, 16'hBD97, 16'hB515, 16'h838E, 16'hBD96, 16'hEEDB, 16'hC596, 16'hFFDF, 16'hF75D, 16'hC514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hE65A, 16'hDE18, 16'hD596, 16'hD5D7, 16'hCD55, 16'hFF1D, 16'hEE1A, 16'hEE19, 16'hE619, 16'hD556, 16'hC4D4, 16'hC515, 16'hC4D4, 16'hC4D4, 16'hCD15, 16'h9B4E, 16'hC4D4, 16'hCD56, 16'hD556, 16'h9B4E, 16'hB451, 16'hFEDC, 16'hF6DD, 16'hFEDC, 16'hC492, 16'hAB4D, 16'hC410, 16'hD514, 16'hCC93, 16'h9B0B, 16'h8248, 16'h7A48, 16'h5985, 16'h4040, 16'h5904, 16'h50C2, 16'h5904, 16'h8249, 16'hABCE, 16'hD514, 16'hF69A, 16'hFF9E, 16'hFF9E, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hD556, 16'hE618, 16'hFF5E, 16'hDD97, 16'h89C6, 16'h8A08, 16'h8A07, 16'h7986, 16'h7185, 16'h6984, 16'h9B4D, 16'hCD14, 16'hBC91, 16'h934C, 16'h6A48, 16'h5986, 16'h5185, 16'h59C6, 16'h59C6, 16'h5185, 16'h4103, 16'h4944, 16'h4944, 16'h5185, 16'h5185, 16'h59C6, 16'h5185, 16'h38C2, 16'h4102, 16'h61C6, 16'h8A89, 16'hB3CF, 16'hEE5A, 16'hFF9F, 16'hFF9F, 16'hC493, 16'hBB8E, 16'hCCD3, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD16, 16'hCCD4, 16'h7A48, 16'hBC92, 16'hD596, 16'h8249, 16'hB492, 16'hCD96, 16'hB492, 16'h5985, 16'h830C, 16'h8B4D, 16'h9C10, 16'hBD14, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hBCD4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB515, 16'h9C11, 16'hA452, 16'hB4D4, 16'h93CF, 16'hAC92, 16'h838E, 16'hB515, 16'hB515, 16'hACD4, 16'hBD56, 16'hBD56, 16'h7B8E,
        16'hAD14, 16'hF75D, 16'hC556, 16'hFF9E, 16'hFFDF, 16'hBCD4, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hDE18, 16'hDDD7, 16'hDDD8, 16'hD5D7, 16'hCD55, 16'hFF1D, 16'hEE1A, 16'hEE19,
        16'hE619, 16'hD597, 16'hC4D4, 16'hC515, 16'hC4D4, 16'hC494, 16'hCD15, 16'h9B4D, 16'hBC93, 16'hD557, 16'hD515, 16'h8ACB, 16'hDD55, 16'hFF1D, 16'hF6DC, 16'hE5D7, 16'hC451, 16'hC451, 16'hD4D3, 16'hABCF, 16'h6103, 16'h6186, 16'h38C3, 16'h2800, 16'h4903, 16'h5185, 16'h4103, 16'h5144, 16'h4903, 16'h3881, 16'h4880, 16'h6102, 16'hAB4C, 16'hDD96, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hF71D, 16'hFFDF, 16'hFF5D, 16'hB38E, 16'h9186, 16'h9A49, 16'h9248, 16'h7985, 16'h8248, 16'hC4D2, 16'hDD96, 16'hBC91, 16'h7248, 16'h4944, 16'h5185, 16'h6207, 16'h7249, 16'h59C6, 16'h5986, 16'h5986, 16'h6A07, 16'h6A48, 16'h59C6, 16'h5185, 16'h5184, 16'h5985, 16'h4903, 16'h4903, 16'h4944, 16'h38C2, 16'h4944,
        16'h8289, 16'hB3CF, 16'hE5D7, 16'hFF9F, 16'hBC92, 16'hBBCF, 16'hD514, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD15, 16'h828A, 16'hB452, 16'hDD97, 16'h828A, 16'hAC51, 16'hCD56, 16'hCD55, 16'h7ACB, 16'h7249, 16'h8B4C, 16'h9C10, 16'hBD14, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hBCD4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hBD15, 16'hA452, 16'h9C10, 16'hB514, 16'h93CF, 16'hAC93, 16'h8B8E, 16'hB4D4, 16'hB515, 16'hACD4, 16'hB556, 16'hBD56, 16'h7B8E, 16'hA4D3, 16'hFFDF, 16'hD5D7, 16'hEF1C, 16'hFFDF, 16'hCD55, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hE659, 16'hCD14, 16'hEE5A, 16'hCD96, 16'hCD14, 16'hFEDD, 16'hEE5A, 16'hEE1A, 16'hE619, 16'hD556, 16'hC4D4, 16'hC515, 16'hC4D4, 16'hC494, 16'hCD16, 16'h934D, 16'hB452, 16'hDD97, 16'hCCD4, 16'h92CB, 16'hEE19, 16'hFF1D, 16'hEE19, 16'hE619, 16'hF6DB, 16'hDD55, 16'h930C, 16'h6A48, 16'h4103, 16'h30C2, 16'h4104, 16'h5144, 16'h4903, 16'h5103, 16'h5103, 16'h61C6, 16'h61C6, 16'h5985, 16'h61C6, 16'h59C6, 16'h5103, 16'h7944, 16'hCC92, 16'hFF1D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hC451, 16'hAB0C, 16'hC3CF, 16'hAACB, 16'h89C6, 16'h928A, 16'hD514, 16'hE5D6, 16'hCCD3, 16'h7A89, 16'h40C2, 16'h6A08, 16'h7ACA, 16'h7ACA, 16'h7289, 16'h6A48, 16'h7A89, 16'h82CB, 16'h7A89, 16'h6A07, 16'h7A89, 16'h7248, 16'h5144, 16'h6A07, 16'h9B8C, 16'h7A48, 16'h5143, 16'h4143, 16'h4143, 16'h4903, 16'h5902, 16'h8A89, 16'hDD97, 16'hBC51, 16'hB3CF, 16'hD4D4, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD516, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD15, 16'h8ACB, 16'hA3D0, 16'hD556, 16'h828A, 16'hA411, 16'hCD56, 16'hCD56, 16'hAC51, 16'h5945, 16'h6A48, 16'h9C0F, 16'hBD14, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB515,
        16'hB4D3, 16'h93D0, 16'hBD15, 16'h9410, 16'hA452, 16'h93CF, 16'hA493, 16'hB556, 16'hA4D4, 16'hB515, 16'hBD96, 16'h83CF, 16'h9C91, 16'hFF9F, 16'hE65A, 16'hDE59, 16'hFFDF, 16'hD618, 16'hDE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9A, 16'hC491, 16'hF71D, 16'hD5D7, 16'hCD55, 16'hFEDC, 16'hEE5A, 16'hEE1A, 16'hEE19, 16'hD556, 16'hC515, 16'hC515, 16'hC4D4, 16'hBC93, 16'hCD56, 16'h9B4E, 16'hB451, 16'hDD97, 16'hBC52, 16'hA38E, 16'hFEDC, 16'hF71D, 16'hF71D, 16'hFF9F, 16'hFF5E, 16'hCD55, 16'h61C5, 16'h30C2, 16'h30C3, 16'h4104, 16'h40C2, 16'h3800, 16'h61C6, 16'h7289, 16'h8B4C, 16'h6207, 16'h5144, 16'h5986, 16'h61C6, 16'h4944, 16'h5144, 16'h4944, 16'h8207, 16'hC451, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65A, 16'hCC52, 16'hF61A, 16'hE516, 16'hA28A, 16'h8A89, 16'hD554, 16'hDDD7, 16'hD554, 16'h8B0B, 16'h3840, 16'h7A8A, 16'h830B, 16'h82CA, 16'h82CA, 16'h7249, 16'h82CA, 16'h7A89,
        16'h82CB, 16'h828A, 16'h7A8A, 16'h8ACB, 16'h82CA, 16'h7249, 16'h5144, 16'hA38D, 16'hCCD2, 16'h9B4C, 16'h5943, 16'h5185, 16'h5144, 16'h4944, 16'h5985, 16'h71C6, 16'h8A49, 16'hC451, 16'hCC93, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD516, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD15, 16'h930C, 16'hA38F, 16'hDD56, 16'h8ACA, 16'hAC51, 16'hCD56, 16'hC555, 16'hC514, 16'h728A, 16'h5145, 16'h8B8D, 16'hBD14, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB515, 16'hB4D4, 16'h93D0, 16'hB4D4, 16'h9C51, 16'hA451, 16'h9410, 16'h9C51, 16'hB556, 16'hA493, 16'hAD15, 16'hBD97, 16'h8C11, 16'h8C10, 16'hF79E, 16'hF71C, 16'hCD96, 16'hFFDF, 16'hE6DB, 16'hC555, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hAB8E, 16'hFF9F, 16'hD596, 16'hD596, 16'hF6DC, 16'hEE5A, 16'hEE5A, 16'hE61A, 16'hCD56, 16'hC515, 16'hC515, 16'hC4D5, 16'hBC93, 16'hCD15, 16'h9B8F, 16'hAC10, 16'hE597, 16'hA38E, 16'hBC92, 16'hFF1D, 16'hF71D, 16'hFF9E, 16'hFF5E, 16'hE618, 16'h6A07, 16'h30C2, 16'h3103, 16'h3903, 16'h2800, 16'h6207, 16'hA40F, 16'hB4D2, 16'hC513, 16'h9BCE, 16'h4943, 16'h6207, 16'h51C6, 16'h59C6, 16'h5185,
        16'h4944, 16'h38C1, 16'h5185, 16'h7206, 16'hBC0F, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'hFF1E, 16'hFE5B, 16'hC3D1, 16'h924A, 16'hD554, 16'hDE17, 16'hDDD6, 16'hBC91, 16'h48C3, 16'h6A08, 16'h82CA, 16'h82CA, 16'h8B0B, 16'h7289, 16'h7A8A, 16'h82CB, 16'h82CA, 16'h7249, 16'h7A8A, 16'h8B0C, 16'h7A8A, 16'h82CB, 16'h8B0B, 16'h6A48, 16'h61C6, 16'hCCD3, 16'hD554, 16'hA3CE, 16'h5944, 16'h6A07, 16'h5185, 16'h6185, 16'h69C6, 16'h4800, 16'h930C, 16'hBC10, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'h930D, 16'hA3CF, 16'hDD96, 16'h828A, 16'hB492, 16'hCD56, 16'hC515, 16'hCD55, 16'hA3CF,
        16'h2800, 16'h7B0B, 16'hB514, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB515, 16'h9C10, 16'hAC93, 16'hA452, 16'h9C51, 16'h9C51, 16'h9410, 16'hB556, 16'hA4D3, 16'hAD15, 16'hBD97, 16'h9452, 16'h8BCF, 16'hEF1D, 16'hFF9E, 16'hC555, 16'hFF9F, 16'hF75D, 16'hBD14, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65A, 16'hA38E, 16'hFF9F, 16'hC555, 16'hD596, 16'hF6DC, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hCD56, 16'hC515, 16'hC515, 16'hC4D5, 16'hBC93, 16'hCD15, 16'hA38F, 16'hA3CF, 16'hDD55, 16'h928A, 16'hDD96, 16'hFF1D, 16'hF75E, 16'hF71D, 16'hD555, 16'h8B0B, 16'h4104, 16'h3103, 16'h3903, 16'h3800, 16'h830B, 16'hC554, 16'hCD95, 16'hC595, 16'hB492, 16'h48C2, 16'h61C6, 16'h6A48, 16'h6A48, 16'h7249, 16'h7249, 16'h6A07, 16'h5184, 16'h61C6, 16'h7248, 16'h7185, 16'hC410, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hF65B, 16'hD492, 16'hCCD3, 16'hE618,
        16'hDDD7, 16'hDDD7, 16'h934D, 16'h48C3, 16'h7ACA, 16'h7A8A, 16'h8B0C, 16'h8B0B, 16'h7A49, 16'h8ACB, 16'h828A, 16'h828A, 16'h8ACB, 16'h8B0C, 16'h82CB, 16'h7249, 16'h82CA, 16'h8B0B, 16'h82CB, 16'h48C2, 16'hA40F, 16'hD595, 16'hCD54, 16'hA3CE, 16'h69C5, 16'h61C6, 16'h4903, 16'h7207, 16'h6145, 16'h79C7, 16'h8208, 16'hC493, 16'hDD56, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD516, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD15, 16'hCD56, 16'h9B4E, 16'hA38E, 16'hD555, 16'h7A49, 16'hBCD3, 16'hCD55, 16'hC515, 16'hC555, 16'hB492, 16'h48C2, 16'h6A8A, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hBD15, 16'hA452, 16'hA452, 16'hAC93, 16'h93CF, 16'hAC93, 16'h93D0, 16'hB555, 16'hA4D4, 16'hACD4, 16'hBD97, 16'h9C93, 16'h83CF, 16'hE6DC, 16'hFFDF, 16'hCD96, 16'hEF1C, 16'hFFDF, 16'hBD14, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC596, 16'hA38D, 16'hFF9E, 16'hAC51, 16'hD5D8, 16'hFF1D, 16'hEE5A, 16'hEE5A, 16'hEE19, 16'hCD56, 16'hC515, 16'hC515, 16'hC515, 16'hBC53, 16'hCD15, 16'hABD0, 16'hA3CF, 16'hBC52, 16'h8207, 16'hEE18, 16'hFF5E, 16'hF6DC, 16'hD514, 16'h7A47, 16'h1800, 16'h2882, 16'h5185, 16'h48C1,
        16'h8B4C, 16'hCD95, 16'hCD95, 16'hC595, 16'hC554, 16'h7ACA, 16'h50C2, 16'h7248, 16'h6A48, 16'h7249, 16'h7A89, 16'h7A89, 16'h7249, 16'h7A89, 16'h6A07, 16'h69C6, 16'h7A48, 16'hB30C, 16'hD514, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hF65B, 16'hEDD8, 16'hF69A, 16'hE5D8, 16'hDDD7, 16'hD595, 16'h6A07, 16'h7249, 16'h8B0C, 16'h82CB, 16'h930C, 16'h7A8A, 16'h82CA, 16'h8ACB, 16'h82CB, 16'h8ACB, 16'h930C, 16'h8ACB, 16'h8ACB, 16'h828A, 16'h82CB, 16'h828A, 16'h930C, 16'h7289, 16'h7ACA, 16'hCD55, 16'hCD95, 16'hCD55, 16'h9B8D, 16'h5944, 16'h6186, 16'h5944, 16'h6145, 16'hB3CF, 16'hC451, 16'hB410, 16'hD515, 16'hD557, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD16,
        16'hCD16, 16'hCD16, 16'hCD56, 16'hA38F, 16'h934D, 16'hC4D3, 16'h7208, 16'hC4D4, 16'hCD55, 16'hC515, 16'hC555, 16'hBCD4, 16'h6A08, 16'h51C7, 16'hACD3, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB515, 16'hAC93, 16'h9C11, 16'hB4D4, 16'h8B8F, 16'hB4D4, 16'h8B8F, 16'hB515, 16'hACD4, 16'hA4D4, 16'hBD56, 16'hA4D4, 16'h83CF, 16'hD659, 16'hFFDF, 16'hD618, 16'hDE99, 16'hFFDF, 16'hC555, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD54, 16'hC451, 16'hFF1D, 16'hAC51, 16'hD5D8, 16'hFF1D, 16'hEE5A, 16'hEE5A, 16'hE619, 16'hCD56, 16'hC515, 16'hC515, 16'hCD15, 16'hBC52, 16'hC515, 16'hB412, 16'h9B4D, 16'h82CB, 16'h8ACA, 16'hF69A, 16'hFF1D, 16'hE618, 16'hB410, 16'h3902, 16'h3944, 16'h4985, 16'h4902, 16'h834C, 16'hCD95, 16'hC595, 16'hC595, 16'hCDD5, 16'hB4D1, 16'h5102, 16'h7207, 16'h7A89, 16'h7248, 16'h7A8A, 16'h7A89, 16'h7A8A, 16'h82CB, 16'h7A8A, 16'h828A, 16'h7208, 16'h6185, 16'hA2CB, 16'hE596, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFEDD, 16'hFEDD, 16'hFEDC, 16'hF65B, 16'hE618, 16'hC514, 16'h6986, 16'h82CB, 16'h82CB, 16'h82CA, 16'h7249, 16'h7A8A, 16'h82CB, 16'h8ACB, 16'h930C, 16'h930C, 16'h8ACB, 16'h828A, 16'h82CB, 16'h82CB, 16'h8B0B, 16'h934D, 16'h9B4D, 16'h82CA, 16'h7A89, 16'hCD54, 16'hCD96, 16'hCD95, 16'hC513, 16'h8A89, 16'h69C6, 16'h6986, 16'h6144, 16'hB3CF, 16'hD493, 16'hDD56, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD56, 16'hABD0, 16'h930C, 16'hBC92, 16'h7249, 16'hC514, 16'hC555, 16'hC515, 16'hC515, 16'hC514, 16'h82CB, 16'h3881, 16'hA451, 16'hB514, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB515, 16'hB4D4, 16'h93D0, 16'hACD3, 16'h8B8E, 16'hB4D4, 16'h93CF, 16'hACD4, 16'hAD15, 16'hA4D4, 16'hBD96, 16'hACD4, 16'h7B8E, 16'hC5D7, 16'hFFDF, 16'hE6DB, 16'hCD96, 16'hFFDF, 16'hD618, 16'hDE59,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hCD14, 16'hDD55, 16'hEEDC, 16'hB4D3, 16'hD5D7, 16'hFF1D, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hCD56, 16'hC515, 16'hC515, 16'hC515, 16'hBC93, 16'hC515, 16'hB452,
        16'h7A89, 16'h48C3, 16'hA38E, 16'hFEDC, 16'hF6DC, 16'hDD96, 16'h38C0, 16'h30C2, 16'h4985, 16'h5185, 16'h59C6, 16'hBD54, 16'hCDD6, 16'hC595, 16'hC595, 16'hC595, 16'h9BCE, 16'h5040, 16'h7A89, 16'h7A89, 16'h7A89, 16'h82CA, 16'h7A89, 16'h82CA, 16'h82CB, 16'h8ACB, 16'h7A8A, 16'h7A48, 16'h7A49, 16'h68C2, 16'hBBCF, 16'hFF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hFEDD, 16'hFEDD, 16'hFEDD, 16'hFEDB, 16'hC4D3, 16'h6144, 16'h82CB, 16'h9BCF, 16'hB4D3, 16'h9BCF, 16'h82CB, 16'h8B0C, 16'h930C, 16'h930C, 16'h8ACC, 16'h8ACB, 16'h8B0C, 16'h8ACB, 16'h934D, 16'h9B8E, 16'h9B4D, 16'h930C, 16'h8ACB, 16'h69C6, 16'hBCD2, 16'hD5D6, 16'hCD95, 16'hCD55, 16'h9B4C, 16'h58C2, 16'h928A, 16'h8207, 16'h9B0D, 16'hCC93, 16'hD515,
        16'hD557, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD15, 16'hAC10, 16'h930C, 16'hB451, 16'h7249, 16'hC514, 16'hC555, 16'hC555, 16'hC515, 16'hC514, 16'h8B0D, 16'h40C1, 16'h9C10, 16'hB515, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D5, 16'h9411, 16'hAC93, 16'h8B8F, 16'hACD4, 16'h9410, 16'hA493, 16'hAD15, 16'hA493, 16'hB556, 16'hAD15, 16'h7B8E, 16'hC597, 16'hFF9E, 16'hF79E, 16'hC556, 16'hFFDF, 16'hE69A, 16'hCD97, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hD5D7, 16'hDDD7, 16'hE659, 16'h9BCF, 16'hD597, 16'hFF1D, 16'hEE5A, 16'hEE5A, 16'hEE19, 16'hCD15, 16'hC515, 16'hC515, 16'hC515, 16'hBC93, 16'hC4D5, 16'hBC93, 16'h828A, 16'h50C2, 16'hB410, 16'hFF1D, 16'hE659, 16'h7248, 16'h1000, 16'h4944, 16'h6A07, 16'h4080, 16'h93CD, 16'hCDD6, 16'hC595, 16'hCD95, 16'hC595, 16'hC595, 16'h82CA, 16'h5903, 16'h7248, 16'h6A07, 16'h7289, 16'h82CA, 16'h82CA, 16'h82CB, 16'h82CA, 16'h82CB, 16'h8ACB, 16'h828A, 16'h8ACB, 16'h7A08, 16'h9248, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hBCD3, 16'h5881, 16'h8B4E, 16'h9C11, 16'hCD97, 16'hCD97, 16'h9BD0, 16'h934D, 16'h934E, 16'h930D, 16'h8ACC, 16'h8B0C, 16'h930C, 16'h934D, 16'h9B8E, 16'h9B4D, 16'h930C, 16'h9B4D, 16'h9B4D, 16'h4800, 16'hAC50, 16'hD5D6, 16'hCD96, 16'hD596, 16'hB40F, 16'h6984, 16'hAB4D, 16'hA2CB, 16'hB3D0, 16'hD4D4, 16'hD515, 16'hDD57, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD16, 16'hCD15, 16'hCD15, 16'hAC11, 16'h930B, 16'hABCF, 16'h830C, 16'hC515, 16'hC555, 16'hC555, 16'hC515, 16'hC514, 16'h8B0D, 16'h59C6, 16'h93CF, 16'hB514, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB515, 16'h9C11, 16'hA452, 16'h9410, 16'hACD4, 16'h9C51, 16'hA492,
        16'hB516, 16'h9C93, 16'hB556, 16'hB515, 16'h838E, 16'hB555, 16'hF79E, 16'hFFDF, 16'hCD96, 16'hF79E, 16'hF75D, 16'hC515, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE18, 16'hF71C, 16'hCD55, 16'hEE5A, 16'h934E,
        16'hD597, 16'hFF1D, 16'hEE1A, 16'hEE5A, 16'hE619, 16'hCD15, 16'hC515, 16'hC515, 16'hC515, 16'hBC93, 16'hC494, 16'hC4D4, 16'h8ACB, 16'h6185, 16'hB410, 16'hFE9B, 16'hA3CE, 16'h000, 16'h51C6, 16'h6A48, 16'h5145, 16'h5944, 16'hBD12, 16'hCDD6, 16'hC5D5, 16'hC5D6, 16'hC5D6, 16'hBD54, 16'h7288, 16'h6A07, 16'h7ACA, 16'h8B8E, 16'h834C, 16'h7A8A, 16'h8ACB, 16'h8B0B, 16'h82CA, 16'h82CA, 16'h930B, 16'h930B, 16'h930C, 16'h9B0C, 16'h7081, 16'hC4D3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC513, 16'h71C7, 16'h9BD0, 16'h93D0, 16'h93D0, 16'h93D1, 16'h9BD0, 16'h938E, 16'h9B8F, 16'h934E, 16'h934D, 16'h934D, 16'h930D, 16'h9B8E, 16'h930D, 16'h930D, 16'h9B4E, 16'h9B8E, 16'h930C,
        16'h6944, 16'hAC50, 16'hD5D6, 16'hD596, 16'hDDD7, 16'hC491, 16'h6984, 16'hB34E, 16'hA2CB, 16'hD4D4, 16'hDD15, 16'hD4D5, 16'hD557, 16'hD556, 16'hD557, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD15, 16'hAC11, 16'h8ACA, 16'hA38E, 16'h82CB, 16'hC515, 16'hC555, 16'hC555, 16'hC555, 16'hC515, 16'h934E, 16'h6A07, 16'h834D, 16'hB514, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB515, 16'hA493, 16'h9C51, 16'h9410, 16'hACD3, 16'hAC93, 16'h8C10, 16'hB556, 16'h9C92, 16'hB555, 16'hB556, 16'h83CF, 16'hAD14, 16'hF75D, 16'hFFDF, 16'hDE19, 16'hEF1C, 16'hFFDF, 16'hC514, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD5D6, 16'hF71C, 16'hC4D2, 16'hEE5A, 16'h9B8E, 16'hD556, 16'hFF1D, 16'hEE5A, 16'hEE5A, 16'hE5D9, 16'hCD15, 16'hC515, 16'hC515, 16'hCD15, 16'hC4D4, 16'hBC93, 16'hCCD5, 16'h930C, 16'h7A07, 16'hB38D, 16'hD4D2, 16'h4903, 16'h59C6, 16'h934B, 16'h7A49, 16'h5144, 16'h7289, 16'hC595, 16'hCDD6, 16'hC5D6, 16'hC5D6, 16'hCDD6, 16'hBD54, 16'h6A07, 16'h7248, 16'h93CF, 16'hEF1C, 16'hCDD8, 16'h728A, 16'h82CB, 16'h934C, 16'h930C, 16'h930C, 16'h9B0C, 16'h9B0C, 16'hA34D, 16'hAB4E, 16'h92CB, 16'h9249,
        16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC555, 16'h71C7, 16'h9C11, 16'hA453, 16'hAC53, 16'hA453, 16'hAC52, 16'h9C11, 16'h9BD0, 16'h934E, 16'h7A89, 16'h934D, 16'h9B8E, 16'h934D, 16'h9B4E, 16'hA38F, 16'h9B8E, 16'h9B4E, 16'hA34D, 16'h7185, 16'hA40F, 16'hD5D6, 16'hCD95, 16'hD5D6, 16'hBC50, 16'h8207, 16'hB34D, 16'hAB0C, 16'hD4D4, 16'hDD15, 16'hD4D5, 16'hD557, 16'hD556, 16'hD557, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD15, 16'hAC11, 16'h8A8A, 16'h930C, 16'h8B0C, 16'hC555, 16'hC515, 16'hC555, 16'hBD14, 16'hC515, 16'h934E, 16'h6A07, 16'h834D, 16'hB514, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4,
        16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB515, 16'hAC93, 16'h9410, 16'h9C51, 16'h9C52, 16'hB514, 16'h838F, 16'hB515, 16'h9C92, 16'hB515, 16'hB556, 16'h8C10, 16'hA4D3, 16'hEF5D, 16'hFFDF, 16'hE69A, 16'hD618, 16'hFFDF, 16'hC555, 16'hEF1B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hDE18, 16'hFF5D, 16'hD514, 16'hE65A, 16'h930C, 16'hCD15, 16'hFF1D, 16'hF65B, 16'hF65B, 16'hE5D8, 16'hC515, 16'hC515, 16'hC515, 16'hCD15, 16'hC4D4, 16'hBC93, 16'hCD15, 16'h9B0D, 16'h71C6, 16'hB38E, 16'h8249, 16'h3902, 16'hABCE, 16'hABCE, 16'h5185, 16'h5985, 16'h838C, 16'hCDD6, 16'hC5D6, 16'hC5D6, 16'hC5D6, 16'hCDD6, 16'hBD13, 16'h6A06, 16'h7248, 16'h834C, 16'hBD55, 16'hA492, 16'h8B4D, 16'h934D, 16'h8B0B, 16'h930B, 16'h9B0C, 16'hA30D, 16'hAB0D, 16'hAB4D, 16'hB38E, 16'hA34E, 16'h8103, 16'hDDD8, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD5D7, 16'h7145, 16'hAC53, 16'hA453, 16'hA494, 16'hAC93, 16'hB494,
        16'hB4D4, 16'hA452, 16'h9BCF, 16'h7289, 16'h8B0C, 16'hA38F, 16'hA38F, 16'hA3D0, 16'h9B8F, 16'h9B4D, 16'hA34E, 16'hA38E, 16'h7185, 16'hC513, 16'hFF5D, 16'hEEDB, 16'hDDD7, 16'hBC0F, 16'h8A07, 16'hCC51, 16'hAB0D, 16'hD4D4, 16'hDD16, 16'hD4D5, 16'hD557, 16'hD556, 16'hD557, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD15, 16'hAC11, 16'h8248, 16'h71C7, 16'hA410, 16'hCD55, 16'hC515, 16'hC515, 16'hBD15, 16'hC515, 16'h938E, 16'h7ACA, 16'h72CB, 16'hACD4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hACD4, 16'hACD4, 16'hB4D4, 16'hB4D4, 16'h9410, 16'h9C11, 16'h9411, 16'hB515, 16'h838E, 16'hACD4, 16'h9C92, 16'hAD15, 16'hB556, 16'h8C11, 16'h9C92, 16'hEF1C, 16'hFFDF, 16'hF75D, 16'hCD96, 16'hFFDF, 16'hD618, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE659, 16'hEEDB, 16'hF69A, 16'hDD55, 16'hEE9A, 16'hA3CF, 16'hCCD4, 16'hFEDD, 16'hF69C, 16'hF65B, 16'hE5D8, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D4, 16'hBC53, 16'hCD15, 16'h930D, 16'h7186, 16'h7A07, 16'h4103, 16'h8ACB, 16'hCC50, 16'h9B0B, 16'h5985, 16'h6144, 16'h9C0F, 16'hCE16, 16'hC5D6, 16'hC5D6, 16'hCDD6, 16'hD5D7, 16'hD5D6, 16'h7248, 16'h7ACA, 16'h938E, 16'h830C,
        16'h830C, 16'h9BCF, 16'hA3D0, 16'h938E, 16'h82CB, 16'h8A8A, 16'hAB4E, 16'hB34E, 16'hB38E, 16'hB38F, 16'hB38F, 16'h9A4A, 16'hBC51, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9A, 16'h81C6, 16'hAC53, 16'hB4D5, 16'hB4D5, 16'hB4D5, 16'hB4D5, 16'hB4D4, 16'hAC94, 16'hA452, 16'h9C11, 16'h938F, 16'hA412, 16'hB452, 16'hAC11, 16'hA3D0, 16'hA3CF, 16'hABCF, 16'hB3CF, 16'h7143, 16'hCD96, 16'hFFDF, 16'hFFDF, 16'hFF5D, 16'hC491, 16'h9A4A, 16'hE4D4, 16'hB34D, 16'hD4D4, 16'hDD16, 16'hD515, 16'hD557, 16'hD556, 16'hD557, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD15, 16'hAC11, 16'h6986, 16'h5945, 16'hB451, 16'hCD55,
        16'hC555, 16'hC515, 16'hBD15, 16'hC515, 16'h938F, 16'h6A48, 16'h6A8A, 16'hACD3, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB515, 16'h93D0, 16'h9410, 16'h8BCF, 16'hB555, 16'h8BD0, 16'hA493, 16'h9451, 16'hAD15, 16'hB556, 16'h8C11, 16'h9411, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hCD97, 16'hFF9E, 16'hEEDB, 16'hD618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD5D7, 16'hF75D, 16'hEE59, 16'hDD96, 16'hD597, 16'hABD0, 16'hD514, 16'hF6DC, 16'hF69C, 16'hF65B, 16'hDDD8, 16'hC4D5, 16'hC515, 16'hC515, 16'hC515, 16'hCD15, 16'hBC52, 16'hCCD5, 16'h9B4E, 16'h48C2, 16'h4944, 16'h69C5, 16'hDD56, 16'hE597, 16'h9ACA, 16'h930B, 16'h8A89, 16'h9BCE, 16'hCE16, 16'hC5D6, 16'hCDD6, 16'hE658, 16'hEEDB, 16'hF71B, 16'h8B4D, 16'h6207, 16'h9410, 16'h9411, 16'h9C11, 16'hA411, 16'h9BD0, 16'hA410, 16'h9BCF, 16'h82CB, 16'hA34D, 16'hB38E, 16'hB38E, 16'hB38F, 16'hB3D0, 16'hAB4E, 16'hAB4E, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h9B4D, 16'hAC11, 16'hBD16, 16'hBD16, 16'hB516, 16'hB4D6, 16'hBD16, 16'hC557, 16'hBD16, 16'hBD16, 16'hB4D5, 16'hBCD5, 16'hBCD5, 16'hAC93, 16'hAC52, 16'hB494, 16'hBC94, 16'hAC11, 16'h7986, 16'hE699, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hA34D, 16'hC410, 16'hF597, 16'hA2CB, 16'hD4D5, 16'hDD16, 16'hD515, 16'hDD57, 16'hD557, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD15, 16'hAC11, 16'h5904, 16'h5986, 16'hBCD3, 16'hC555, 16'hC555, 16'hC555, 16'hBD15, 16'hC515, 16'h830C, 16'h7ACB, 16'h72CA, 16'hA492, 16'hB4D5, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB515, 16'h9C11, 16'h9410, 16'h8BD0, 16'hB555, 16'h8BD0, 16'h9C92, 16'h9411, 16'hAD14, 16'hB556, 16'h8C51, 16'h8BCF, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hDE18, 16'hF71C, 16'hF75D, 16'hCD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hE659, 16'hF71D, 16'hEEDB, 16'hE618, 16'hCD14, 16'hAC11, 16'hE5D8, 16'hEE9B, 16'hF6DC, 16'hF65B, 16'hDD98, 16'hC4D5, 16'hC515, 16'hC515, 16'hC515, 16'hCD15, 16'hBC93, 16'hC4D4, 16'h7A8A, 16'h38C2, 16'h51C6, 16'hA34D, 16'hEE19, 16'hFF1D, 16'hDD97, 16'hAB4B,
        16'h9ACB, 16'h9B4C, 16'hCDD6, 16'hC596, 16'hE69A, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hB4D3, 16'h5983, 16'h9C51, 16'h9411, 16'hA453, 16'hA453, 16'hA453, 16'hA452, 16'hA411, 16'hA3D0, 16'h8B0C, 16'hA38F, 16'hB3D0, 16'hB3CF, 16'hBC11, 16'hBB90, 16'hA28B, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD55, 16'h9B4E, 16'hCD98, 16'hC557, 16'hC558, 16'hC557, 16'hC557, 16'hCD58, 16'hC558, 16'hCD58, 16'hCD57, 16'hC557, 16'hC517, 16'hCD98, 16'hCD98, 16'hBD16, 16'hB494, 16'h9B4F, 16'hA38E, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hE619, 16'hBB4D, 16'hEE19, 16'hED98, 16'h9A8A, 16'hDD15, 16'hDD56, 16'hD515, 16'hDD57, 16'hD557, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556,
        16'hCD56, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD15, 16'hB451, 16'h5040, 16'h7A8A, 16'hC555, 16'hC555, 16'hC555, 16'hC515, 16'hBD15, 16'hC514, 16'h7ACC, 16'h830C, 16'h830C, 16'hA492, 16'hB4D5, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hACD4, 16'hB515, 16'hA493, 16'h8BD0, 16'h838E, 16'hAD15, 16'h9411, 16'h9C52, 16'h9411, 16'hAD14, 16'hB556, 16'h9452, 16'h838E, 16'hCDD8, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hDE59, 16'hFF9E, 16'hCD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9A, 16'hEEDB, 16'hEEDB, 16'hFF5E, 16'hE618, 16'hC515, 16'hAC50, 16'hEE59, 16'hEE5A, 16'hF6DC, 16'hF65B, 16'hDD97, 16'hC4D5, 16'hC515, 16'hC515, 16'hC515, 16'hCD15, 16'hBC93, 16'hC4D4, 16'hAC10, 16'h4103, 16'h5185, 16'h7A48, 16'hD514, 16'hFEDC, 16'hFEDD, 16'hC451, 16'hAB0B, 16'hAB4D, 16'hC514, 16'hEE9A, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'h6142, 16'hA452, 16'h9C53, 16'hA453, 16'hA494, 16'hA494, 16'hA453, 16'hA453, 16'hB494, 16'hAC12, 16'hA412, 16'hB453, 16'hBC94, 16'hBC53, 16'hBC52, 16'hAACB, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hA38D, 16'hCD57, 16'hDDDA, 16'hD5D9, 16'hD5D9, 16'hD5D9, 16'hD5D9, 16'hD5D9, 16'hD5D9, 16'hD599, 16'hCD99, 16'hCD98, 16'hEE9C, 16'hFF5F, 16'hF71E, 16'hE65B, 16'hCD57, 16'hDE19, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD4D4, 16'hED97, 16'hFF1D, 16'hE597, 16'hA2CC, 16'hDD57, 16'hDD56, 16'hD515, 16'hDD57, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD16, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD56, 16'hCD15, 16'hCD15, 16'hB452, 16'h3000, 16'h938F, 16'hCD56, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hB4D3, 16'h59C7, 16'h7ACB, 16'h7B0B, 16'h9C52, 16'hB4D5, 16'hACD4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB514, 16'hB514, 16'hACD5, 16'hB515, 16'hACD3, 16'h8BD0, 16'h838E, 16'hAD15, 16'h9C52, 16'h9451, 16'h9C92, 16'hA4D4, 16'hB556, 16'h9C93, 16'h83CF, 16'hBD96, 16'hFFDF,
        16'hFFDF, 16'hEF1C, 16'hCDD7, 16'hFFDF, 16'hC555, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE58, 16'hF71C, 16'hEEDC, 16'hFFDF, 16'hE618, 16'hBC92, 16'hAC51, 16'hEE5A, 16'hE5D8, 16'hFEDD, 16'hF65B, 16'hDD97, 16'hC4D5, 16'hC515, 16'hC515,
        16'hC515, 16'hCD15, 16'hBC93, 16'hAC11, 16'h82CC, 16'h5186, 16'h51C7, 16'h5184, 16'h930A, 16'hDD96, 16'hFF1E, 16'hEE5A, 16'hBBCF, 16'hAB4C, 16'hD555, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h8B4C, 16'h8B8F, 16'hACD5, 16'hAD16, 16'hB4D6, 16'hB4D6, 16'hACD5, 16'hB4D5, 16'hB4D5, 16'hC557, 16'hC517, 16'hC557, 16'hCD98, 16'hCD57, 16'hDE1A, 16'hDD97, 16'hEE9B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD595, 16'hBC52, 16'hE61A, 16'hDE1A, 16'hDE1A, 16'hDE1A, 16'hDE1A, 16'hDE1A, 16'hDE1A, 16'hDDDA, 16'hDDDA, 16'hD5DA, 16'hD5DA, 16'hDE1B, 16'hE65C, 16'hE65C, 16'hFE9D, 16'hFF1D, 16'hFFDF, 16'hFF9F, 16'hF65B, 16'hED56, 16'hEDD7, 16'hFEDC, 16'hE597,
        16'hB34D, 16'hE557, 16'hDD56, 16'hD515, 16'hDD57, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD16, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD56, 16'hCD15, 16'hCD15, 16'hAC11, 16'h5945, 16'hB493, 16'hC555, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hA451, 16'h6208, 16'h7B0C, 16'h72CA, 16'h9C11, 16'hB4D5, 16'hACD4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hACD4, 16'hB514, 16'hAD15, 16'hACD5, 16'hB4D5, 16'hACD4, 16'h9410, 16'h8BCF, 16'hAD14, 16'hA4D3, 16'h9411, 16'h9C93, 16'hA4D4, 16'hB556, 16'hA4D4, 16'h8C10, 16'hB514, 16'hF79E, 16'hFFDF, 16'hFF9E, 16'hCDD7, 16'hFFDF, 16'hCD97, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hE659, 16'hF71C, 16'hF71D, 16'hFFDF, 16'hE618, 16'hB411, 16'hA410, 16'hEE9B, 16'hDD97, 16'hFEDC, 16'hF65B, 16'hD597, 16'hC4D5, 16'hC515, 16'hC515, 16'hC515, 16'hCD15, 16'hC4D4, 16'hB452, 16'hAC51, 16'h51C7, 16'h9C92, 16'h5A8A, 16'h4901, 16'hABCE, 16'hF65A, 16'hFEDD, 16'hF69B, 16'hC451, 16'hC451, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD617, 16'h7A89, 16'hACD5, 16'hAD16, 16'hBD17, 16'hC557, 16'hC557, 16'hBD17, 16'hC558, 16'hD599, 16'hD599, 16'hCD99, 16'hD599, 16'hD5D9, 16'hDE5B, 16'hDDD9, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hD556, 16'hD598, 16'hE65B, 16'hDE1A, 16'hDE1A, 16'hDE1A, 16'hDE1A, 16'hDE1A, 16'hDE1A, 16'hDE1A, 16'hDE1A, 16'hDE1A, 16'hD5DA, 16'hE61A, 16'hCC94, 16'hDCD5, 16'hFF9E, 16'hFF9F, 16'hF69C, 16'hF61A, 16'hFE5A, 16'hF65A, 16'hFEDD, 16'hE556, 16'hAB0D, 16'hE557, 16'hDD56, 16'hD515, 16'hDD57, 16'hD557, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD56, 16'hCD15, 16'hCD15, 16'hAC11, 16'h7A8A, 16'hC514, 16'hC515, 16'hC515, 16'hC515, 16'hC514, 16'hC515, 16'h9BD0, 16'h6A09, 16'h830C, 16'h830C, 16'h9410, 16'hB515, 16'hACD4, 16'hACD4, 16'hB514, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hAD15, 16'hAD15, 16'hAD15, 16'hAD15,
        16'h9411, 16'h838E, 16'h9C93, 16'hAD14, 16'h8BD0, 16'h9C93, 16'hA493, 16'hB556, 16'hA4D4, 16'h83CF, 16'hA492, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hCD96, 16'hF75D, 16'hDE59, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hE69A, 16'hEEDB, 16'hFF5E,
        16'hFFDF, 16'hE619, 16'hB411, 16'hA410, 16'hF6DC, 16'hD556, 16'hF6DC, 16'hF65B, 16'hD597, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D4, 16'hB452, 16'hBCD4, 16'h5186, 16'hAD14, 16'h8C11, 16'h2800, 16'h59C4, 16'hC492, 16'hFE9B, 16'hFEDD, 16'hF69B, 16'hE658, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hA40E, 16'h9C11, 16'hBD57, 16'hBD16, 16'hC558, 16'hC598, 16'hCD98, 16'hD5D9, 16'hD5D9, 16'hD5DA, 16'hD61A, 16'hDE1A, 16'hDE1A, 16'hDE1A, 16'hD557, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hD597, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B,
        16'hEE5C, 16'hE598, 16'hC34F, 16'hF69B, 16'hFFDF, 16'hFEDC, 16'hFE5B, 16'hF65B, 16'hF65B, 16'hFEDC, 16'hFF1D, 16'hDD15, 16'hB34D, 16'hE557, 16'hDD56, 16'hD515, 16'hDD57, 16'hD557, 16'hD557, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD56, 16'hCD15, 16'hCD15, 16'hB451, 16'h7A49, 16'hBCD4, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'h8B4D, 16'h7ACB, 16'h830C, 16'h8B4D, 16'h8BCF, 16'hB515, 16'hACD4, 16'hAD15, 16'hB514, 16'hB4D4, 16'hAD14, 16'hAD14, 16'hAD14, 16'hAD14, 16'hAD15, 16'hAD15, 16'hB515, 16'h9C52, 16'h838E, 16'h9C93, 16'hB556, 16'h83CF, 16'h9C93, 16'hA493, 16'hAD15, 16'hAD15, 16'h8C11, 16'h9C51, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'hE6DB, 16'hE6DB, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE659, 16'hF71C, 16'hEE9A, 16'hFF9E, 16'hFFDF, 16'hE65A, 16'hABD0, 16'hAC51, 16'hFF5D, 16'hD556, 16'hF69C, 16'hF65B, 16'hD557, 16'hC4D5, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D5, 16'hB412, 16'hBCD4, 16'h59C7, 16'hA4D3, 16'h9C93, 16'h5208, 16'h59C7, 16'h8A8A, 16'hE597, 16'hFEDC, 16'hFF1D, 16'hF6DC, 16'hEE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE699, 16'h7A89, 16'hBD57, 16'hC598, 16'hC558, 16'hCD98, 16'hD5D9, 16'hDE1A, 16'hDE1A, 16'hDE5B,
        16'hDE5B, 16'hE65B, 16'hE69B, 16'hE65B, 16'hDDD9, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hE65C, 16'hEE1B, 16'hDD16, 16'hCBD2, 16'hEE5A, 16'hFF5E, 16'hF69B, 16'hED97, 16'hED97, 16'hED98, 16'hFE9B, 16'hFEDC, 16'hFEDD, 16'hD4D4, 16'hB38E, 16'hE598, 16'hDD57, 16'hDD16, 16'hDD57, 16'hD557, 16'hD557, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD15, 16'hCD15, 16'hB452, 16'h7A8A, 16'hBCD4, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hBCD4, 16'h728A, 16'h830C, 16'h82CC, 16'h8B4D, 16'h838F,
        16'hAD15, 16'hACD4, 16'hAD15, 16'hACD4, 16'hACD4, 16'hACD5, 16'hAD15, 16'hACD4, 16'hACD4, 16'hACD5, 16'hACD5, 16'hAD15, 16'h9C93, 16'h838E, 16'h9C92, 16'hB556, 16'h8BD0, 16'h9C93, 16'hA4D4, 16'hAD15, 16'hAD15, 16'h9452, 16'h9410, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'hDE59, 16'hEEDB, 16'hD5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hDE18, 16'hF75D, 16'hE699, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'h92CB, 16'hAC92, 16'hFF9E, 16'hCD56, 16'hF65B, 16'hF69B, 16'hD557, 16'hC4D5, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hB452, 16'hBCD4, 16'h728A, 16'h9C92, 16'h9C92, 16'h734D, 16'h6ACA, 16'h5902, 16'hBC10, 16'hF65A, 16'hFF1D, 16'hEE1A, 16'hEE19, 16'hFF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC554, 16'h9B8E, 16'hD5D9, 16'hDE1A, 16'hDE1A, 16'hE65B, 16'hE65B, 16'hE69C, 16'hE69C, 16'hE69C, 16'hE69C, 16'hEE9C, 16'hE65B, 16'hE69B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hEEDC, 16'hEE9C, 16'hEE5C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE5B, 16'hF69C, 16'hEE1A, 16'hDCD4, 16'hF5D8, 16'hFE9C, 16'hF65B, 16'hF65A, 16'hED98, 16'hEDD8, 16'hEDD8, 16'hF65A, 16'hFF1D, 16'hFEDD, 16'hCC52, 16'hBBD0, 16'hE598, 16'hDD57, 16'hD515, 16'hDD57, 16'hD557, 16'hD557, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD15, 16'hCD15, 16'hCD15, 16'hB411, 16'h7A8A, 16'hC514, 16'hC515, 16'hC515, 16'hC515, 16'hC555, 16'hA451, 16'h6A49, 16'h9C10, 16'h8B4D, 16'h938E, 16'h8BCF, 16'hAD15, 16'hACD4, 16'hAD15, 16'hACD4, 16'hACD4, 16'hACD4, 16'hACD4, 16'hACD4, 16'hAD15, 16'hACD5, 16'hACD5, 16'hAD15, 16'hA4D4, 16'h7B4E, 16'h9411, 16'hB557, 16'h8C10, 16'h9C93, 16'h9C93, 16'hAD15, 16'hA4D5, 16'h8C11, 16'hA492, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hD618, 16'hEF1C, 16'hC596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hE69A, 16'hEEDC, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'h9ACC, 16'hA411, 16'hFF9F, 16'hD596, 16'hEE1A, 16'hF69B, 16'hD557, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hCD15, 16'hB452, 16'hC4D4, 16'h7ACB, 16'h8C10, 16'hAD14, 16'h7B8E, 16'h7B8E, 16'h5903, 16'h8248, 16'hDD55, 16'hFEDD, 16'hFF1D, 16'hFEDD, 16'hF69B, 16'hFEDC, 16'hFF5E, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD554, 16'hBC12, 16'hE65B, 16'hEE9C, 16'hE69C, 16'hE69C, 16'hE69C, 16'hE69C, 16'hEE9C, 16'hEEDC, 16'hEE9C, 16'hEEDC, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF69B, 16'hFF1D, 16'hEE5B, 16'hF69C, 16'hEE5A, 16'hE557, 16'hED98, 16'hEDD9, 16'hE516, 16'hFF1D, 16'hF61A, 16'hDCD4, 16'hE4D5, 16'hEE19, 16'hFEDC, 16'hFEDC, 16'hFEDD, 16'hFEDD, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hBC11, 16'hBC11, 16'hE598, 16'hDD57, 16'hD4D5, 16'hD556, 16'hD557, 16'hD557, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD15, 16'hCD15, 16'hC515, 16'hAC11,
        16'h82CA, 16'hC514, 16'hC515, 16'hC515, 16'hC515, 16'hC555, 16'h834D, 16'h72CB, 16'hAC93, 16'h7ACB, 16'h8B4D, 16'h838E, 16'hAD15, 16'hACD4, 16'hAD15, 16'hACD4, 16'hACD4, 16'hACD4, 16'hACD4, 16'hACD5, 16'hAD15, 16'hAD15, 16'hAD15, 16'hAD15, 16'hACD4, 16'h838E, 16'h9452, 16'hBD97, 16'h9452, 16'h9C92, 16'h9C93, 16'hAD15, 16'hA4D5, 16'h8C12, 16'hB514, 16'hCD96, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD5D8, 16'hEF1C, 16'hCD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hF71C, 16'hE69A, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h92CC, 16'hB4D3, 16'hFFDF, 16'hCD96, 16'hE619, 16'hF65B, 16'hD556, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hBC53, 16'hBC93, 16'h8B4D, 16'h7B8E, 16'hAD15, 16'h7B8E, 16'h9CD3, 16'h6249, 16'h5902, 16'hAB8D, 16'hFE9B, 16'hFEDC, 16'hFE9C, 16'hFE9B, 16'hFE9B, 16'hFE9C, 16'hFF1D, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE5D7, 16'hCCD4, 16'hDDD9, 16'hE65C, 16'hE69C, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hF65A, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF6DC, 16'hF65A, 16'hF69C, 16'hFEDC, 16'hEE19, 16'hFF1D, 16'hFF1D, 16'hF69C, 16'hF65A, 16'hFEDC, 16'hFF1D, 16'hFF1D, 16'hFEDC, 16'hFEDD, 16'hFEDD, 16'hFF1D, 16'hFEDC, 16'hB38F, 16'hC452, 16'hE598, 16'hE597, 16'hD4D4, 16'hD516, 16'hDD57, 16'hD557, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC515, 16'hA410, 16'h82CB, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hB4D3, 16'h4185, 16'h838E, 16'hB4D4, 16'h7ACB, 16'h834D, 16'h838E, 16'hAD15, 16'hACD4, 16'hAD15, 16'hACD5, 16'hACD4, 16'hACD4, 16'hACD4, 16'hAD15, 16'hAD15, 16'hAD15, 16'hAD15, 16'hAD15, 16'hAD15, 16'h83CF, 16'h8C11, 16'hBD97, 16'h9452, 16'h9452, 16'hA4D4, 16'hAD15, 16'hAD15, 16'h8C11, 16'hC597, 16'hD5D7, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hD618, 16'hEF1C, 16'hD5D7, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'hF75D, 16'hDDD8, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h8ACB, 16'hB4D3, 16'hFFDF, 16'hD5D7, 16'hDD97, 16'hF65B, 16'hCD56, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hBC94, 16'hC493, 16'h938E, 16'h7B4E, 16'hB556,
        16'h7B8F, 16'hA4D4, 16'h8BD0, 16'h4902, 16'h7184, 16'hD514, 16'hFE9B, 16'hF6DC, 16'hF65B, 16'hF5D9, 16'hF65A, 16'hFE5B, 16'hFE9C, 16'hFF1D, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'hDDD7, 16'hDD56, 16'hEE9B, 16'hEE9C, 16'hE65B, 16'hDDD9, 16'hE69B, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF6DC, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFEDC, 16'hFEDC, 16'hFEDD, 16'hFF1D, 16'hFEDC, 16'hFEDD, 16'hFF1D, 16'hF65A, 16'hB34E, 16'hCC53, 16'hE598, 16'hDD97, 16'hD4D4, 16'hD515, 16'hD557, 16'hD556, 16'hD556,
        16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD15, 16'hCD15, 16'hC515, 16'hC515, 16'hA410, 16'h82CB, 16'hC515, 16'hC515, 16'hBD14, 16'hC515, 16'h9C10, 16'h2800, 16'h9C51, 16'hB4D4, 16'h7B0B, 16'h834D, 16'h838F, 16'hAD15, 16'hACD4, 16'hAD15, 16'hAD15, 16'hACD4, 16'hACD5, 16'hAD15, 16'hAD15, 16'hAD15, 16'hAD15, 16'hAD15, 16'hAD15, 16'hAD15, 16'h8BD0, 16'h83D0, 16'hBD97, 16'h9C93, 16'h8C11, 16'h9C93, 16'hA4D4, 16'hAD15, 16'h8410, 16'hCE18, 16'hD618, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hD5D8, 16'hE6DB, 16'hC555, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hE69A, 16'hFF9E, 16'hDDD8, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h828B, 16'hAC92, 16'hFFDF, 16'hDE19, 16'hD515, 16'hF65A, 16'hCD56, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hBC94, 16'hBC53, 16'h9BD0, 16'h6ACB, 16'hB555, 16'h734E, 16'h9C93, 16'hAD15, 16'h6249, 16'h5903, 16'hA30C, 16'hF65A, 16'hFF1D, 16'hF619, 16'hED57, 16'hF5D8, 16'hDCD4, 16'hF598, 16'hF61A, 16'hFEDC, 16'hFF5E, 16'hFF5D, 16'hEE9A, 16'hFF5E, 16'hFF5D, 16'hF69A, 16'hFF1D, 16'hEE5B, 16'hE619, 16'hF6DC, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1D, 16'hFEDC, 16'hFF1D, 16'hF6DC, 16'hFF1D, 16'hFEDC, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFEDC, 16'hFEDC, 16'hF69B, 16'hFF1D, 16'hF6DB, 16'hFEDC, 16'hFEDD, 16'hFEDD, 16'hED97, 16'hBB4E, 16'hD493, 16'hE598, 16'hDD97, 16'hD4D5, 16'hD515, 16'hD557, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD56, 16'hCD15, 16'hCD15, 16'hC515, 16'hC515, 16'hAC11, 16'h7ACB, 16'hC515, 16'hBD15, 16'hBD14, 16'hBD14, 16'h6ACB, 16'h5A49, 16'hACD3, 16'hACD4, 16'h7B0C, 16'h834D, 16'h838E, 16'hAD15, 16'hACD4, 16'hAD15, 16'hAD15, 16'hACD5, 16'hACD5, 16'hAD15, 16'hAD15, 16'hAD15, 16'hAD15, 16'hAD15, 16'hAD15, 16'hB515, 16'h9411, 16'h83CF, 16'hB597, 16'hA4D4, 16'h9452, 16'h9CD4, 16'hA514,
        16'hAD55, 16'h7BCF, 16'hCE19, 16'hE69A, 16'hCDD7, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'hDE5A, 16'hC555, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hEEDB, 16'hF71D, 16'hDE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h828A, 16'hA492, 16'hFFDF, 16'hE69A, 16'hCD15, 16'hEE1A,
        16'hCD56, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC4D5, 16'hBC53, 16'h9BD0, 16'h7B0C, 16'hB555, 16'h7BCF, 16'h9C93, 16'hB556, 16'h8C10, 16'h3840, 16'h8207, 16'hEDD8, 16'hF69B, 16'hF65B, 16'hFE5B, 16'hED97, 16'hE555, 16'hF597, 16'hED56, 16'hFE9B, 16'hFF5E, 16'hF69B, 16'hEE19, 16'hFF1D, 16'hFF1D, 16'hF69B, 16'hFF5D, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF65A, 16'hF619, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5D, 16'hFF1D, 16'hFF1D, 16'hFEDC, 16'hFF1D, 16'hFEDC, 16'hF6DC, 16'hFF1D, 16'hFF1D, 16'hFEDC, 16'hFEDC, 16'hF69B, 16'hFEDC, 16'hFEDB, 16'hF69B, 16'hFF1D,
        16'hFEDC, 16'hF65B, 16'hE516, 16'hBB4E, 16'hD493, 16'hE598, 16'hDD97, 16'hD4D4, 16'hD515, 16'hD597, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD15, 16'hC515, 16'hC515, 16'hA3D0, 16'h8B0C, 16'hC555, 16'hBD14, 16'hBD15, 16'h9C10, 16'h2000, 16'h8BD0, 16'hAD15, 16'hACD4, 16'h7B0C, 16'h8B8E, 16'h838F, 16'hAD15, 16'hACD5, 16'hA515, 16'hA515, 16'hACD4, 16'hACD5, 16'hA515, 16'hAD15, 16'hAD15, 16'hACD5, 16'hACD5, 16'hAD15, 16'hAD16, 16'h9C52, 16'h7B4E, 16'hB557, 16'hA4D4, 16'h9452, 16'h9C93, 16'hA4D4, 16'hAD56, 16'h83D0, 16'hCE19, 16'hF75D, 16'hC554, 16'hFFDF, 16'hFFDF, 16'hE69B, 16'hD618, 16'hCD96, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE18, 16'hFF5E, 16'hE6DB, 16'hE65A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h828A, 16'hAC52, 16'hFFDF, 16'hF71C, 16'hCD15, 16'hE5D9, 16'hCD56, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hB452, 16'hA411, 16'h6A8A, 16'hB555, 16'h8410, 16'h9452, 16'hB556, 16'hACD4, 16'h6B0C, 16'h4800, 16'hB411, 16'hFE9B, 16'hF69B, 16'hFEDC, 16'hFEDC, 16'hF65A, 16'hF65A, 16'hF65A, 16'hFF1D, 16'hFF1D, 16'hFEDD, 16'hFEDD, 16'hF71D, 16'hFF5D, 16'hFF5D, 16'hFF5D, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF65A, 16'hED57, 16'hFF1D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1C, 16'hFF1D, 16'hF6DC, 16'hFF1D, 16'hFEDD, 16'hF69B, 16'hFF1D, 16'hFF1D, 16'hFEDC, 16'hF69B, 16'hF69B, 16'hF69B, 16'hFEDC, 16'hF65A, 16'hFF1D, 16'hFEDC, 16'hF69B, 16'hFE9B, 16'hD4D4, 16'hC38F, 16'hD4D4, 16'hE598, 16'hDD98, 16'hD4D4, 16'hD515, 16'hD557, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD15, 16'hCD15, 16'hC4D4, 16'hC515, 16'h9BD0, 16'h8B0C, 16'hC515, 16'hBD15, 16'hAC92, 16'h3904, 16'h6ACB, 16'hACD4, 16'hA4D4, 16'hACD4, 16'h7B0C, 16'h7B0D, 16'h838F, 16'hAD15, 16'hACD5, 16'hA515, 16'hA515, 16'hACD4, 16'hACD4, 16'hA515, 16'hAD15,
        16'hAD15, 16'hACD5, 16'hACD5, 16'hAD15, 16'hAD16, 16'h9C93, 16'h7B4F, 16'hB556, 16'hAD15, 16'h8C11, 16'h9C93, 16'h9CD4, 16'hB556, 16'h83D0, 16'hC5D7, 16'hFF9F, 16'hC554, 16'hFF9E, 16'hFFDF, 16'hEF1C, 16'hD5D7, 16'hC555, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD5D7, 16'hFFDF,
        16'hDE19, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'h8249, 16'hB492, 16'hFFDF, 16'hF75D, 16'hCD15, 16'hE5D9, 16'hCD56, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hB453, 16'hAC11, 16'h728A, 16'hAD15, 16'h9492, 16'h8C10, 16'hB556, 16'hB515, 16'h9C52, 16'h4080, 16'h9B0C, 16'hF5D9, 16'hF65B, 16'hFEDD, 16'hEE5A, 16'hF65A, 16'hF69B, 16'hFEDC, 16'hFF1D, 16'hF6DC, 16'hF69B, 16'hF6DC, 16'hFF1D, 16'hFF5D, 16'hFF1D, 16'hFF5D, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hF69B, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF1D, 16'hFF1C, 16'hFF1C, 16'hF6DC, 16'hFF1D,
        16'hF69B, 16'hFF1D, 16'hFF1D, 16'hF69B, 16'hF69B, 16'hF65B, 16'hF65A, 16'hFEDC, 16'hF65A, 16'hFF1D, 16'hFF1C, 16'hF69A, 16'hFEDC, 16'hFE9B, 16'hD452, 16'hC390, 16'hD4D5, 16'hE598, 16'hDD98, 16'hD4D4, 16'hD515, 16'hD557, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD16, 16'hC515, 16'hBCD4, 16'hBCD5, 16'hA411, 16'h830C, 16'hBD14, 16'hB4D3, 16'h5A49, 16'h3904, 16'h9C92, 16'hACD4, 16'hA4D4, 16'hACD4, 16'h730C, 16'h7B4D, 16'h838F, 16'hAD15, 16'hACD5, 16'hA515, 16'hA515, 16'hACD5, 16'hACD5, 16'hA515, 16'hA4D5, 16'hA515, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hAD15, 16'hA4D4, 16'h7B8F, 16'hB556, 16'hAD16, 16'h8C11, 16'h9C93, 16'h9493, 16'hAD56, 16'h83D0, 16'hBD97, 16'hFFDF, 16'hCD96, 16'hEF1C, 16'hFFDF, 16'hF75D, 16'hCD97, 16'hCD95, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hDE59, 16'hFFDF, 16'hDE18, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'h8249, 16'hB493, 16'hFF9E, 16'hFF5E, 16'hCD15, 16'hDD98, 16'hCD56, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hBC93, 16'hB452, 16'h728A, 16'hA4D3, 16'h9493, 16'h8410, 16'hB556, 16'hAD15, 16'hA4D4, 16'h628A, 16'h7185, 16'hE556, 16'hFE9C, 16'hF619, 16'hF69B, 16'hF69B, 16'hF65A, 16'hFF1D, 16'hFEDC, 16'hF69A, 16'hF69B, 16'hFF1C, 16'hFF1D, 16'hFEDC,
        16'hFF1C, 16'hFF1D, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF1D, 16'hF71C, 16'hFF1C, 16'hF6DC, 16'hFF1D, 16'hF69B, 16'hFF1D, 16'hFF1D, 16'hF69B, 16'hF69B, 16'hF65A, 16'hF619, 16'hFE9B, 16'hF65A, 16'hF6DC, 16'hFF1D, 16'hF65A, 16'hFEDC, 16'hFF1D, 16'hF619, 16'hD452, 16'hCBD1, 16'hD4D5, 16'hE598, 16'hDD98, 16'hD4D5, 16'hCD15, 16'hD557, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD16, 16'hCD16, 16'hCD16, 16'hC515, 16'hC515, 16'hBCD4, 16'hBD15, 16'h9BD0, 16'h834C, 16'hB4D3, 16'h6A8A, 16'h2800, 16'h9C51, 16'hAD15, 16'hA4D4, 16'hACD4,
        16'hACD4, 16'h730C, 16'h834D, 16'h8BCF, 16'hAD15, 16'hAD15, 16'hAD15, 16'hA515, 16'hACD5, 16'hACD5, 16'hA515, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hAD15, 16'hA4D4, 16'h7B8F, 16'hAD56, 16'hAD56, 16'h8C11, 16'h9C93, 16'h9452, 16'hAD56, 16'h7B8F, 16'hC5D7, 16'hFFDF, 16'hDE18, 16'hDE59, 16'hFFDF, 16'hF79E, 16'hC555, 16'hCD55, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65A, 16'hEF1C, 16'hFF9E, 16'hD596, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h9B8E, 16'hBCD2, 16'hF75D, 16'hFF9F, 16'hD597, 16'hD557, 16'hCD56, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hBC94, 16'hB492, 16'h72CB, 16'h9C51, 16'hA514, 16'h83CF, 16'hB556, 16'hAD15, 16'hB556, 16'h8BCF, 16'h5000, 16'hD4D4, 16'hF619, 16'hF65A, 16'hFE9B, 16'hF65A, 16'hFEDD, 16'hFEDC, 16'hF69A, 16'hF69B, 16'hF69B, 16'hFF1D, 16'hF6DC, 16'hFEDC, 16'hFF1D, 16'hFF1D, 16'hFF5D, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF1D, 16'hFEDC, 16'hFF1D, 16'hFEDC, 16'hFF1D, 16'hF69B, 16'hFEDD, 16'hFF1E, 16'hF69B, 16'hF69B, 16'hF69B, 16'hF65A, 16'hF69B, 16'hFE9C, 16'hF69B, 16'hFF1D, 16'hF69B, 16'hFEDC, 16'hFEDD, 16'hF69B, 16'hEDD9, 16'hDC52, 16'hD452, 16'hDD15, 16'hDD97, 16'hDD98, 16'hD515, 16'hCD15, 16'hD557, 16'hD556, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD16, 16'hC516, 16'hC516, 16'hC515, 16'hBCD4, 16'hBCD4, 16'h9BCF, 16'h7B0C, 16'h5A48, 16'h3904, 16'h9411, 16'hAD15, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D4, 16'h730C, 16'h7B0C, 16'h8BD0, 16'hAD15, 16'hAD15, 16'hAD15, 16'hA515, 16'hAD15, 16'hAD15, 16'hA515, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hAD15, 16'hA4D5, 16'h838F, 16'hAD16, 16'hAD56, 16'h8C11, 16'h9492, 16'h9452, 16'hB597, 16'h7B8F, 16'hC5D8, 16'hFFDF, 16'hE6DB, 16'hD5D7, 16'hFFDF, 16'hFF9F, 16'hC555, 16'hAC51, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD618, 16'hFF9F, 16'hF71D, 16'hD5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'hA410, 16'hC514, 16'hEEDC, 16'hFFDF, 16'hDDD8, 16'hCD16, 16'hCD16, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hBCD4, 16'hB493, 16'h8B4D, 16'h9410, 16'h9CD3, 16'h738E, 16'hB556, 16'hAD16, 16'hAD15, 16'h8BD0, 16'h61C6, 16'hAB4D,
        16'hF5D8, 16'hF65A, 16'hEE19, 16'hFEDC, 16'hFEDD, 16'hF61A, 16'hF65A, 16'hF65A, 16'hFF1D, 16'hF6DC, 16'hF6DB, 16'hFF1D, 16'hF71C, 16'hFF5D, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF5D, 16'hF71C, 16'hFF1D, 16'hFF1C, 16'hFF1D, 16'hF69B, 16'hFEDC, 16'hFF5E, 16'hF6DC, 16'hF69B, 16'hF69B, 16'hF65A, 16'hF69B, 16'hFF1D, 16'hF65B, 16'hFF1D, 16'hF69B, 16'hFEDC, 16'hFF1D, 16'hF65B, 16'hF6DC, 16'hEDD9, 16'hD452, 16'hCBD0, 16'hDD15, 16'hDD97, 16'hDD97, 16'hCCD5, 16'hCCD4, 16'hD597, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC516, 16'hC516, 16'hC515,
        16'hC4D5, 16'hBCD4, 16'hBCD4, 16'h9BCF, 16'h1000, 16'h5208, 16'hA493, 16'hAD15, 16'hA4D4, 16'hA515, 16'hA4D5, 16'hA4D5, 16'hA4D4, 16'h734D, 16'h7B4C, 16'h8BD0, 16'hAD16, 16'hAD15, 16'hAD15, 16'hA515, 16'hAD15, 16'hAD15, 16'hA515, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA515, 16'hAD15, 16'h83D0, 16'hA515, 16'hB597, 16'h8C11, 16'h9493, 16'h9452, 16'hB556, 16'h7B8F, 16'hD659, 16'hFFDF, 16'hF75D, 16'hCD96, 16'hFFDF, 16'hFFDF, 16'hD5D7, 16'hAC0F, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hE65A, 16'hFFDF, 16'hEE9B, 16'hE659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCDD7, 16'hB4D3, 16'hC555, 16'hE659, 16'hFFDF, 16'hE619, 16'hCD15, 16'hCD16, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hBCD4, 16'hAC52, 16'h9BCF, 16'h838E, 16'hA4D3, 16'h7BCF, 16'hAD15, 16'hAD16, 16'hAD15, 16'h9C52, 16'h61C6, 16'h92CC, 16'hFE9C, 16'hEDD9, 16'hF69B, 16'hFF1D, 16'hF61A, 16'hF65A, 16'hF659, 16'hFEDC, 16'hF6DC, 16'hF69B, 16'hFF1D, 16'hF6DC, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF1C, 16'hFF5D, 16'hFF5D, 16'hFF5D, 16'hF6DC, 16'hFEDC, 16'hFF5E, 16'hFF1C, 16'hF6DC, 16'hFF1C, 16'hF65A, 16'hF69B, 16'hFF1D, 16'hFEDC, 16'hF69C, 16'hF6DC, 16'hF6DC, 16'hFF1D, 16'hF69B, 16'hF69C, 16'hFF1D, 16'hEDD8, 16'hDC53, 16'hC411, 16'hDD56, 16'hDD97, 16'hDD97, 16'hCCD5, 16'hC4D4, 16'hD597, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC516, 16'hC515, 16'hC515, 16'hC515, 16'hBCD5, 16'hB4D4, 16'hBD14, 16'h938F, 16'h6249, 16'hACD4, 16'hAD15, 16'hA4D5, 16'hA515, 16'hA4D5, 16'hA4D4, 16'hA4D5, 16'hA4D4, 16'h7B4E, 16'h834D, 16'h8BD0, 16'hAD16, 16'hAD15, 16'hAD15, 16'hA515, 16'hAD15, 16'hAD15, 16'hA515, 16'hA515, 16'hA515, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA515, 16'hAD15, 16'h8BD0, 16'hA515, 16'hB597, 16'h8C52, 16'h9493, 16'h9493, 16'hB556, 16'h734D, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hC555, 16'hF75E, 16'hFFDF,
        16'hD5D7, 16'hBC92, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hEEDB, 16'hFFDF, 16'hD5D7, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCDD7, 16'hB514, 16'hD5D7, 16'hD5D7, 16'hFFDF, 16'hE659, 16'hC4D5, 16'hCD15, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515,
        16'hC515, 16'hB452, 16'hAC11, 16'h6249, 16'h9CD3, 16'h7BCF, 16'hAD15, 16'hAD16, 16'hAD15, 16'h8BD0, 16'h6A8A, 16'h79C7, 16'hE597, 16'hFEDC, 16'hFEDC, 16'hF65A, 16'hF65A, 16'hF61A, 16'hFEDB, 16'hFEDC, 16'hF69B, 16'hFF1D, 16'hF6DC, 16'hFF1C, 16'hFF1D, 16'hFF5D, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5D, 16'hFF5E, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF5D, 16'hFF1D, 16'hFF5D, 16'hF69B, 16'hF6DC, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFEDC, 16'hFF1D, 16'hF6DC, 16'hFEDC, 16'hFF1D, 16'hFF1D, 16'hE597, 16'hDC53, 16'hC411, 16'hDD57, 16'hDD97, 16'hD597, 16'hCD15,
        16'hCCD5, 16'hD557, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC516, 16'hC515, 16'hC515, 16'hC515, 16'hBCD4, 16'hB4D4, 16'hBCD4, 16'h938E, 16'h834D, 16'hAD15, 16'hA4D5, 16'hA4D5, 16'hA515, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D4, 16'h7B8E, 16'h7B0C, 16'h8C11, 16'hAD16, 16'hAD15, 16'hAD15, 16'hA515, 16'hAD15, 16'hAD15, 16'hA515, 16'hA515, 16'hA515, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA515, 16'hAD15, 16'h8BD1, 16'hA515, 16'hB597, 16'h9493, 16'h8C52, 16'h9452, 16'hAD56, 16'h730C, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hD5D7, 16'hEEDB, 16'hFFDF, 16'hD617, 16'hA3CF, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hF75D, 16'hFFDF, 16'hDDD7, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD5D7, 16'hC555, 16'hDE59, 16'hC514, 16'hFFDF, 16'hEE9A, 16'hC4D4, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hB452, 16'hB452, 16'h6A89, 16'h9492, 16'h83CF, 16'hACD4, 16'hAD15, 16'hAD15, 16'hAD15, 16'h9C11, 16'h7800, 16'hDD56, 16'hFF5E, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF69B, 16'hFEDC, 16'hF69B, 16'hFF1D, 16'hFEDC, 16'hF6DC, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5D, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5D, 16'hFF5D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hDD55, 16'hDC94, 16'hC411, 16'hDD97, 16'hD557, 16'hD557, 16'hD515, 16'hCD15, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC556, 16'hC516, 16'hC516, 16'hC516, 16'hC515, 16'hB4D4, 16'hB494, 16'hBCD4, 16'h8B4D, 16'h838F, 16'hAD15, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D4, 16'h7B4D, 16'h730C, 16'h8C11, 16'hAD16, 16'hAD15, 16'hA515, 16'hA515, 16'hAD15, 16'hAD15, 16'hA515, 16'hA515, 16'hA515, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA515, 16'hAD15, 16'h8BD1, 16'hA515,
        16'hB597, 16'h9452, 16'h8C52, 16'h9452, 16'hAD15, 16'h730C, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hDE18, 16'hDE59, 16'hFFDF, 16'hD618, 16'h8B4D, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'hFF9E, 16'hFFDF, 16'hCD96, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD96, 16'hC555, 16'hEEDB,
        16'hC4D3, 16'hFF9F, 16'hEE9B, 16'hC4D4, 16'hC515, 16'hCD16, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hB493, 16'hB452, 16'h830C, 16'h8C10, 16'h8C10, 16'hA4D4, 16'hAD15, 16'hA515, 16'hAD15, 16'h9C11, 16'h6840, 16'hDD56, 16'hFE9B, 16'hF69A, 16'hF65A, 16'hF69B, 16'hFF1C, 16'hF69C, 16'hFF1D, 16'hFF1D, 16'hF6DB, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5D,
        16'hFF5D, 16'hFF5E, 16'hFF5D, 16'hFF5D, 16'hFF1D, 16'hD4D4, 16'hD452, 16'hC412, 16'hDD97, 16'hD557, 16'hD597, 16'hCCD5, 16'hC4D4, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC516, 16'hC515, 16'hC515, 16'hC516, 16'hBD15, 16'hB4D4, 16'hB4D4, 16'hBCD4, 16'h830C, 16'h8BD0, 16'hAD15, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D4, 16'h734D, 16'h6ACB, 16'h9452, 16'hAD16, 16'hA515, 16'hA515, 16'hA515, 16'hAD15, 16'hAD15, 16'hA515, 16'hA515, 16'hA515, 16'hA515, 16'hA515, 16'hA515, 16'hA515, 16'hAD15, 16'h8BD1, 16'hA515, 16'hB597, 16'h8C52, 16'h8C52, 16'h9CD4, 16'hA515, 16'h730C, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hE69B, 16'hD5D7, 16'hFFDF, 16'hDE59, 16'hA451, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hD5D7, 16'hFFDF, 16'hFF9E, 16'hCD55, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD14, 16'hBD14, 16'hEEDC, 16'hB451, 16'hFF9E, 16'hEEDB, 16'hC4D4, 16'hC515, 16'hCD56, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hBCD4, 16'hB452, 16'h938F, 16'h734C, 16'h8C10, 16'h9C93, 16'hAD15, 16'hA4D5, 16'hAD15, 16'hA452, 16'h6840, 16'hCCD3, 16'hFEDC, 16'hF69A, 16'hF69B, 16'hFEDC, 16'hFEDC, 16'hFF1D, 16'hFF5D, 16'hFF1D, 16'hFF1D, 16'hFF5D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5D, 16'hCC52, 16'hCBD0, 16'hC453, 16'hDD98, 16'hD557, 16'hD597, 16'hCCD5, 16'hC4D4, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC516, 16'hC516, 16'hC516, 16'hC515, 16'hC515, 16'hC515, 16'hBCD5, 16'hB4D4, 16'hB4D4, 16'hB514, 16'h7B0C, 16'h8C11, 16'hAD15, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D4, 16'h7B4E, 16'h730C, 16'h9452, 16'hAD16, 16'hA515, 16'hA516, 16'hA516,
        16'hAD15, 16'hAD15, 16'hA515, 16'hA515, 16'hA515, 16'hA515, 16'hA515, 16'hA515, 16'hA515, 16'hA515, 16'h8C11, 16'hA4D5, 16'hB597, 16'h8C11, 16'h8C51, 16'h9493, 16'h9C93, 16'h8BCF, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hC555, 16'hFFDF, 16'hDE59, 16'hB4D3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C,
        16'hE69A, 16'hFFDF, 16'hF75C, 16'hD5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB4D3, 16'hB4D3, 16'hF75D, 16'hB451, 16'hFF5D, 16'hF6DC, 16'hC4D4, 16'hBCD4, 16'hCD16, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hBCD5, 16'hB453, 16'hA410, 16'h6B0B, 16'h9451, 16'h9C93, 16'hAD15, 16'hA515, 16'hA515, 16'hA494, 16'h6945, 16'hBC51, 16'hFEDC, 16'hFEDC, 16'hFF1D, 16'hFEDC, 16'hFF1D, 16'hFF5D, 16'hFF5D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF5D, 16'hD452, 16'hCBD0, 16'hCC93, 16'hDD98, 16'hD557, 16'hD597, 16'hCCD5, 16'hC4D4, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC516, 16'hC516, 16'hC516, 16'hC515, 16'hC515, 16'hC515, 16'hBCD4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'h7B0B, 16'h8C11, 16'hAD15, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'h9CD4, 16'h734D, 16'h730C, 16'h9C93, 16'hAD16, 16'hA515, 16'hA516, 16'hA516, 16'hAD15, 16'hAD15, 16'hA516, 16'hA515, 16'hA515, 16'hA515, 16'hA515, 16'hA515, 16'hA515, 16'hA515, 16'h8C52, 16'hA515, 16'hB598, 16'h8C52, 16'h8C11, 16'h9C93, 16'h9452, 16'hA451, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hBCD3, 16'hFF9E, 16'hDE59, 16'hBD14, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hC618, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hEEDB, 16'hFFDF, 16'hE6DB, 16'hCD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBCD3, 16'hBD14, 16'hFF9E, 16'hB451, 16'hF71C, 16'hF6DC, 16'hC4D4, 16'hBCD4, 16'hCD16, 16'hC515, 16'hC515, 16'hC516, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hB453, 16'hAC52, 16'h628A, 16'h8C10, 16'h9C93, 16'hAD15, 16'hA515, 16'hA515, 16'hACD4, 16'h6A08, 16'hA30C, 16'hFEDB, 16'hFF5E, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E,
        16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF5D, 16'hCC11, 16'hC390, 16'hCCD4, 16'hDD97, 16'hD557, 16'hD557, 16'hCCD5, 16'hC494, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC516, 16'hC516, 16'hC516, 16'hC515, 16'hC515, 16'hBD15, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'h7ACB, 16'h9452, 16'hAD16, 16'hA4D5, 16'hA4D5,
        16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA515, 16'h9C93, 16'h730D, 16'h734D, 16'hA4D4, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hAD15, 16'hAD15, 16'hA516, 16'hA516, 16'hA516, 16'hA515, 16'hA515, 16'hA515, 16'hA516, 16'hA515, 16'h8C11, 16'hA516, 16'hB598, 16'h9452, 16'h83D0, 16'h9493, 16'h8411, 16'hA492, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC555, 16'hEF1C, 16'hD618, 16'hBD14, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h7BCF, 16'h7BCF, 16'hD69A, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'hF75D, 16'hFFDF, 16'hDE59, 16'hD618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDE, 16'hC513, 16'hC515, 16'hFF9F, 16'hB492, 16'hE65A, 16'hF6DC, 16'hBCD3, 16'hB493, 16'hCD16, 16'hC515, 16'hC515, 16'hC516, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hB493, 16'hB493, 16'h72CB, 16'h838E, 16'h9C93, 16'hAD15, 16'hA515, 16'hA515, 16'hAD15, 16'h82CB, 16'h9A8A, 16'hF6DB, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9F, 16'hF71D, 16'hBB8F, 16'hC3D0, 16'hCD15, 16'hD557, 16'hD557, 16'hD557, 16'hCCD5, 16'hC494, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC516, 16'hC516, 16'hC516, 16'hBD16, 16'hBD15, 16'hBD15, 16'hBCD5, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'h6A89, 16'h9C93, 16'hA515, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA515, 16'h9493, 16'h734D, 16'h7B4D, 16'hA4D5, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA515, 16'hAD15, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hAD16, 16'h8C11, 16'hA516, 16'hBDD8, 16'h8C52, 16'h7BCF, 16'h8C52, 16'h9451, 16'hBD55, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCDD7, 16'hE69A, 16'hCDD7, 16'hBD54, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8C51, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD618, 16'hFFDE, 16'hFFDF, 16'hD5D7, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hC514, 16'hC514, 16'hFF9F, 16'hBD14, 16'hDDD8, 16'hF6DC, 16'hC4D4, 16'hAC52, 16'hCD56, 16'hC515, 16'hC516, 16'hC516, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hB493, 16'hB493, 16'h838E, 16'h5A48, 16'h9C92, 16'hAD15,
        16'hA515, 16'hA515, 16'hAD15, 16'h8B4E, 16'h79C6, 16'hEE5A, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF71D, 16'hC3CF, 16'hBB8F, 16'hD515, 16'hD557, 16'hCD56, 16'hD557, 16'hCCD5, 16'hC4D4, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC516, 16'hC516, 16'hBD16, 16'hBD15,
        16'hBD15, 16'hBD15, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hAC93, 16'h6A8A, 16'hA4D4, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA515, 16'h9452, 16'h7B8D, 16'h7BCF, 16'hA515, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA515, 16'hA515, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'h8C11, 16'hAD56, 16'hB598, 16'h8410, 16'h7BCF, 16'h9492, 16'h9C52, 16'hC596, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'hDE19, 16'hC555, 16'hC596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hD596, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hCD14, 16'hC514, 16'hFF9E, 16'hC596, 16'hD596, 16'hF6DC, 16'hC514, 16'hAC52, 16'hCD56, 16'hC515, 16'hC516, 16'hC516, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hBCD4, 16'hAC92, 16'h93CF, 16'h5A07, 16'h9C92, 16'hAD15, 16'hAD15, 16'hA515, 16'hAD16, 16'h9C11, 16'h6880, 16'hD597, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF1D, 16'hC3CF, 16'hB38F, 16'hD556, 16'hD557, 16'hCD56, 16'hCD56, 16'hC4D5, 16'hC4D4, 16'hCD56, 16'hCD56, 16'hC516, 16'hC516, 16'hC516, 16'hBD16, 16'hBD15, 16'hBD15, 16'hBD15, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D5, 16'hAC92, 16'h72CB, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA516, 16'h8C11, 16'h7B8E, 16'h83CF, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA515, 16'hA515, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hAD16, 16'hA516, 16'h8411, 16'hAD56, 16'hB597, 16'h8411, 16'h7BD0, 16'h9492, 16'hA4D3, 16'hCDD6, 16'hFF9E, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hE71B, 16'hCD96, 16'hBD14, 16'hD618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hE65A, 16'hFFDF, 16'hFFDF, 16'hCD55, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hC514, 16'hC514, 16'hF71D, 16'hCDD7, 16'hC514, 16'hF6DB, 16'hC515, 16'hAC52, 16'hCD56, 16'hC516, 16'hC516,
        16'hC516, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hBCD5, 16'hB492, 16'h9C10, 16'h4985, 16'h83CF, 16'hAD15, 16'hAD15, 16'hAD15, 16'hAD16, 16'hA493, 16'h6102, 16'hC4D3, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hAB0C, 16'hAB8F, 16'hD557,
        16'hCD56, 16'hCD56, 16'hCD56, 16'hC4D4, 16'hC4D4, 16'hCD56, 16'hC556, 16'hC516, 16'hC516, 16'hC516, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D5, 16'h9C51, 16'h628A, 16'hA515, 16'hA4D5, 16'hA515, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA516, 16'h8C11, 16'h7B8E, 16'h83D0, 16'hAD16, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA515, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hAD16, 16'hAD16, 16'h8411, 16'hAD97, 16'hB597, 16'h7B8F, 16'h8C11, 16'h8410, 16'hB555, 16'hCDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hC514, 16'hA40F, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hCD55, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hCD55, 16'hD596, 16'hE69B, 16'hDE59, 16'hBC93, 16'hF69B, 16'hCD15, 16'hAC11, 16'hCD56, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hAC52, 16'hB4D3, 16'h6249, 16'h734D, 16'hAD15, 16'hAD15, 16'hAD15, 16'hAD16, 16'hAD15, 16'h8ACB, 16'hA34C, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hEF1C, 16'hD5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5D, 16'hBC10, 16'hDE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'h81C7, 16'hABCF, 16'hD597, 16'hCD56, 16'hCD56, 16'hCD16, 16'hBCD4, 16'hBCD4, 16'hCD56, 16'hC516, 16'hC516, 16'hC516, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBCD5, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB4D5, 16'h9410, 16'h6B0C, 16'hAD16, 16'hA4D5, 16'hA515, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA4D5, 16'hA515, 16'h83D0, 16'h734D, 16'h8C11, 16'hAD16, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hAD16, 16'hAD16,
        16'hAD16, 16'hA516, 16'h8452, 16'hB597, 16'hB557, 16'h7BD0, 16'h8410, 16'h83D0, 16'hC596, 16'hCE17, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAC92, 16'h8ACA, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hCE59, 16'hB596, 16'hA514, 16'h9492, 16'h9492, 16'h8410, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE19, 16'hF75D, 16'hFFDF, 16'hFF9F, 16'hC514, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hEE9B, 16'hDE18, 16'hE659, 16'hE659, 16'hE6DB, 16'hB451, 16'hF69B, 16'hC4D4, 16'h9BCF, 16'hCD16, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hAC52, 16'hB4D3, 16'h834D, 16'h51C7, 16'h9C93, 16'hAD55, 16'hAD15, 16'hAD15, 16'hAD16, 16'h9BD0, 16'h70C0, 16'hE659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'h9148, 16'hCD14, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD5D7, 16'h9248, 16'h9ACB, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'h7185, 16'hAC10, 16'hD557, 16'hCD56, 16'hCD56, 16'hC516, 16'hBCD5, 16'hBCD4, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hB4D4, 16'hB4D4, 16'hACD4, 16'hB515, 16'h838E, 16'h7B4E, 16'hAD16, 16'hA4D5, 16'hA516, 16'hA515, 16'hA515, 16'hA515, 16'hA515, 16'hA515, 16'h83CF, 16'h7B8D, 16'h9493, 16'hAD16, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hAD16, 16'hAD16, 16'hA516, 16'hA516, 16'hA516, 16'hAD16, 16'hAD16, 16'hAD57, 16'hA516, 16'h8C52, 16'hBD98, 16'hA516, 16'h83D0, 16'h6B0D, 16'h9C93, 16'hC555, 16'hD699, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hACD2, 16'h82CB, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h9492, 16'h8410, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h8410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD596, 16'hFF9E, 16'hFFDF, 16'hFF9E, 16'hC4D4, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE659, 16'hD618, 16'hE69A, 16'hD5D7, 16'hF71C, 16'hB451, 16'hEE5A, 16'hCD15, 16'hA3D0, 16'hC515, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hC515, 16'hC515, 16'hC515, 16'hC516, 16'hAC52, 16'hAC51, 16'h9C10, 16'h72CC, 16'h628B, 16'hB555, 16'hAD15, 16'hAD15, 16'hAD16, 16'hACD4, 16'h79C6, 16'hC4D2, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE18, 16'h7945, 16'hA30D, 16'hDE19, 16'hFF5D, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hE69A, 16'hD5D7, 16'hA38E, 16'h8208, 16'hC555, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9A, 16'h5800, 16'hB452, 16'hD557, 16'hCD16, 16'hCD56, 16'hC516, 16'hBCD4, 16'hBCD4, 16'hC516, 16'hC516, 16'hC516, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB515, 16'h7B4C, 16'h83D0, 16'hAD56, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'h9CD4, 16'h7B8E, 16'h7B8E, 16'h9494, 16'hAD17,
        16'hAD16, 16'hAD16, 16'hAD16, 16'hA516, 16'hA516, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD57, 16'hA515, 16'h8C52, 16'hBDD8, 16'hA4D4, 16'h7B8F, 16'h630C, 16'hCE18, 16'hBD55, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD55, 16'h9BCF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hBDD7, 16'hA514, 16'h9CD3, 16'h9CD3, 16'hAD55, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'hB596, 16'hAD55, 16'hBDD7, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h9492, 16'h8C51, 16'h8C51, 16'h8C51, 16'h9492, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFF9E, 16'hD5D7, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hCD15, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE18, 16'hD5D7, 16'hF75D, 16'hCD96, 16'hF75D, 16'hAC51, 16'hEE5A, 16'hD556, 16'hA38F, 16'hC515, 16'hCD56, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hC515, 16'hC515, 16'hC515, 16'hC516, 16'hB493, 16'hAC92, 16'h9C11, 16'h9C52, 16'h628A, 16'h83CF, 16'hB556, 16'hAD16, 16'hAD15, 16'hB516, 16'hA3CF, 16'h8A06, 16'hE618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hCD56, 16'hAB8F, 16'hAB8E, 16'hA38F, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE99, 16'hC514, 16'hC555, 16'hDE59, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAC50, 16'h5000, 16'hBC93, 16'hCD56, 16'hCD16, 16'hCD56, 16'hC516, 16'hBCD4, 16'hBCD4, 16'hC516, 16'hC516, 16'hBD16, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hB4D4, 16'hB4D4, 16'hB4D5, 16'hB514, 16'h6249, 16'h8C11, 16'hAD56, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'h9C94, 16'h7B8E, 16'h7B8E, 16'hA515, 16'hAD16, 16'hA516, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD56, 16'hAD56, 16'hAD56, 16'hAD56, 16'hAD56, 16'hAD57, 16'hAD56, 16'hAD57, 16'h9CD5, 16'h9493, 16'hB598, 16'h9493, 16'h738E, 16'h7BCF, 16'hDE59, 16'hB514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD55, 16'hAC51, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hF79E, 16'hB596, 16'h8C51, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h8410, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h9CD3, 16'h8410, 16'h8C51, 16'h8C51, 16'h8C51, 16'h8410, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h8C51, 16'h9492, 16'h9492, 16'hC618, 16'hE71C, 16'hD69A, 16'h8C51, 16'h8C51, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hDE18, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hBCD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD618, 16'hD618, 16'hFFDF, 16'hCD55, 16'hF75D, 16'hB492, 16'hDDD8, 16'hD596, 16'h9B8E, 16'hC515, 16'hCD56, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hC515, 16'hC516, 16'hBCD5, 16'hA451, 16'hA451, 16'h9C51, 16'hB515, 16'h62CB, 16'h8BD0, 16'hB516, 16'hAD16, 16'hAD16, 16'hB4D4, 16'h8A08, 16'hA38D,
        16'hFF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF75D, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD96, 16'h4800, 16'h6A07, 16'hC4D4, 16'hCD57, 16'hC516, 16'hC516, 16'hC515, 16'hB494, 16'hBCD4, 16'hC516, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hB4D5, 16'hB4D4, 16'hB4D4, 16'hB515, 16'hACD4, 16'h4985, 16'h9412,
        16'hAD56, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hAD16, 16'h9453, 16'h6B0C, 16'h7B8F, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hB557, 16'h9CD5, 16'h9CD4, 16'hB598, 16'hA4D4, 16'h7BCF, 16'h9C93, 16'hC556, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB514, 16'hBD14, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h9492, 16'h8C51, 16'h9492, 16'h8C51, 16'h8C51, 16'h8C51, 16'h8C51, 16'h8410, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'hBDD7, 16'hBDD7, 16'hCE59, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h8C51, 16'h9492, 16'h8C51, 16'h8410, 16'h9492, 16'h9492, 16'h8410, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h9492, 16'hE71C, 16'hFFDF, 16'hFFDF,
        16'hF79E, 16'h9492, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'hDE19, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hBC93, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE17, 16'hDE59, 16'hFFDF, 16'hCD96, 16'hEEDB, 16'hBD14, 16'hCD55, 16'hD596, 16'h9B8F, 16'hC4D4, 16'hCD56, 16'hC556, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hC515, 16'hC515, 16'hA411, 16'hB4D3, 16'h9410, 16'hB556, 16'hAD15, 16'h7B8F, 16'h838F, 16'h9C93, 16'hAD16, 16'hB516, 16'hA3D0, 16'h8185, 16'hD554, 16'hFFDE, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCDD7, 16'h1800, 16'h61C7, 16'h7A8A, 16'hC4D4, 16'hC556, 16'hC556, 16'hC556, 16'hC515, 16'hB4D4, 16'hBCD4, 16'hC516, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hB4D5, 16'hB4D4, 16'hB4D4, 16'hB515, 16'h9C52, 16'h4185, 16'h9C93, 16'hAD16, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hAD56, 16'h8C11, 16'h734D, 16'h83CF, 16'hAD57, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD56, 16'hA516, 16'hAD16, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hB557, 16'h9C94, 16'h9CD5, 16'hB597, 16'hA4D4, 16'h6B4D, 16'hB555, 16'hAC92, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA491, 16'hD618, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h9492, 16'h8410, 16'hA514, 16'hDEDB, 16'hEF5D, 16'hE71C, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hA514, 16'h8410, 16'h8C51, 16'h8C51, 16'h8410, 16'h8C51, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8410, 16'h9492, 16'h8C51, 16'hC618, 16'hDEDB, 16'hA514, 16'h8C51, 16'h8C51, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8C51, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hC4D4, 16'hFFDE, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD5D7, 16'hDE59, 16'hFFDF, 16'hD618, 16'hDE5A, 16'hCD96, 16'hCD14, 16'hD596, 16'hA3CF, 16'hBCD4, 16'hCD56, 16'hC556, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hC515, 16'hCD16,
        16'hA411, 16'hAC92, 16'h93D0, 16'hAD15, 16'hAD16, 16'hB516, 16'hA4D4, 16'hA4D4, 16'hAD16, 16'hAD16, 16'hB515, 16'h8B0D, 16'h7A07, 16'hDDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCDD7, 16'h000, 16'h5208, 16'h93D0, 16'h828B, 16'hC515, 16'hC556, 16'hC556, 16'hC516, 16'hBD15, 16'hB4D4, 16'hBCD4, 16'hC515, 16'hBD15, 16'hBD15,
        16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB515, 16'h8BCF, 16'h51C6, 16'hA4D4, 16'hAD57, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hA516, 16'hAD16, 16'h7B8E, 16'h734D, 16'h8C11, 16'hAD57, 16'hAD16, 16'hAD56, 16'hAD56, 16'hAD56, 16'hA516, 16'hAD16, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hB597, 16'h9493, 16'hA516, 16'hAD56, 16'h83D0, 16'h7BCF, 16'hAD14, 16'hB514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h93CF, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9CD3, 16'h8C51, 16'h9492, 16'h8C51, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hF79E, 16'h9CD3, 16'h9492, 16'h8C51, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hEF5D,
        16'h8C51, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hCE59, 16'h8C51, 16'h8C51, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8C51, 16'h8C51, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hC4D3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD5D7, 16'hDE59, 16'hFFDF, 16'hE69A, 16'hD618, 16'hD5D7, 16'hB452, 16'hD556, 16'hA3CF, 16'hBC93, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hCD56, 16'hAC52, 16'hAC92, 16'h9410, 16'hA4D4, 16'hAD16, 16'hAD15, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD15, 16'hAD16, 16'hACD4, 16'h6A49, 16'h8248, 16'hDE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD54, 16'h000, 16'h5A49, 16'hAD14, 16'h9C51, 16'h828A, 16'hCD16, 16'hC516, 16'hC516, 16'hC516, 16'hBD15, 16'hB493, 16'hBCD5, 16'hC516, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hB4D4, 16'hACD4, 16'hB4D4, 16'hB515, 16'h7B0C, 16'h5207, 16'hA4D4, 16'hAD57, 16'hAD16, 16'hAD16, 16'hAD16, 16'hA516, 16'hAD57, 16'h9C93, 16'h7B8E, 16'h7B8E, 16'h9452, 16'hB557, 16'hAD16, 16'hAD57, 16'hAD57, 16'hAD57, 16'hA516, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hB557, 16'h9493, 16'hB597, 16'h9CD4, 16'h5ACB, 16'h8C51, 16'h838D, 16'hE6DB,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h7248, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8410, 16'h9492, 16'h8C51, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8410, 16'h9492, 16'h8C51, 16'hBDD7, 16'hC618, 16'h9492, 16'h9492, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8C51, 16'h8C51, 16'hDEDB, 16'hFFDF, 16'hCE59, 16'h8C51, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h9492, 16'h8410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65A, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hC4D4, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD5D7, 16'hDE99, 16'hFFDF, 16'hEF1C, 16'hC555, 16'hD5D7, 16'hB492, 16'hD556,
        16'hABCF, 16'hB493, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hCD56, 16'hBCD4, 16'hA451, 16'hA451, 16'h9452, 16'hAD16, 16'hAD16, 16'hAD15, 16'hAD15, 16'hAD16, 16'hAD15, 16'hAD15, 16'hAD16, 16'hACD4, 16'h6A48, 16'h8A8A, 16'hE618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hB4D3, 16'h000, 16'h62CB, 16'hAD14, 16'hAD56,
        16'h8B8F, 16'h8ACB, 16'hC556, 16'hC516, 16'hC516, 16'hC516, 16'hBD15, 16'hAC93, 16'hBCD5, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hB515, 16'hB515, 16'hACD4, 16'hACD4, 16'hB515, 16'hAC93, 16'h6249, 16'h7B0C, 16'hA4D5, 16'hAD57, 16'hAD16, 16'hAD17, 16'hAD57, 16'hAD16, 16'hAD57, 16'h8411, 16'h8410, 16'h734D, 16'hA515, 16'hB557, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD56, 16'hAD16, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hB557, 16'hAD57, 16'h8C53, 16'hB597, 16'h9493, 16'h634D, 16'h738D, 16'hB514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h8248, 16'hE6DA, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h9492, 16'h8C51, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hEF5D, 16'hDEDB, 16'hC618, 16'hB596, 16'hE71C, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hD69A,
        16'h8C51, 16'h9492, 16'h9CD3, 16'hFFDF, 16'hDEDB, 16'h8C51, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8C51, 16'h8C51, 16'hD69A, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h9492, 16'hE71C, 16'hFFDF, 16'hEF5D, 16'hB596, 16'h8C51, 16'h9492, 16'h9492, 16'h9CD3, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hBC93, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD5D7, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hBD14, 16'hDDD7, 16'hBC93, 16'hCD15, 16'hAC10, 16'hB452, 16'hCD16, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC516, 16'hCD16, 16'hC4D5, 16'h9BD0, 16'hAC92, 16'h9411, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD15, 16'hAD15, 16'hAD15, 16'hAD16, 16'hACD4, 16'h7249, 16'h79C5, 16'hDDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'h8B4D, 16'h000, 16'h5A8A, 16'hAD14, 16'hA4D3, 16'hB556, 16'h8B8E, 16'h8B0D, 16'hCD57, 16'hC516, 16'hC556, 16'hBD15, 16'hBCD5, 16'hAC53, 16'hBCD5, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hB515, 16'hB4D5, 16'hB4D4, 16'hB515, 16'h9C11, 16'h72CB, 16'h838E, 16'hA4D5, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD16, 16'h734E, 16'h8C52, 16'h6B0C, 16'hAD56, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD56, 16'hAD16, 16'hAD57, 16'hAD57, 16'hB557, 16'hB557,
        16'hB557, 16'hAD57, 16'hAD57, 16'hB598, 16'hAD16, 16'h9493, 16'hB598, 16'h8411, 16'h5ACB, 16'h7B4C, 16'hEF5C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB513, 16'hA3CE, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hC618, 16'hA514, 16'h9CD3, 16'h8C51, 16'h8410, 16'h8410, 16'h8410, 16'h8C51, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h9492, 16'h8C51, 16'hF79E, 16'hE71C, 16'h8410, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h9492, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h8C51, 16'h9492, 16'h9492, 16'hAD55, 16'h8C51, 16'h8C51, 16'h9492, 16'h8C51, 16'h9492, 16'h7BCF, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE18, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hC4D3, 16'hFF9E,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD5D7, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hCDD7, 16'hCD96, 16'hB452, 16'hCD15, 16'hB411, 16'hAC11, 16'hC515, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC516, 16'hCD16, 16'h9BD0, 16'hAC92, 16'h93D0, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD15, 16'hACD5, 16'hAD15, 16'hAD15, 16'hAD16, 16'hACD4, 16'h6A49, 16'h6103, 16'hD596, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hCD96, 16'h5185, 16'h000, 16'h20C1, 16'h8C91, 16'hAD55, 16'h9452, 16'hBD97, 16'h8C10, 16'h934E, 16'hCD57, 16'hC516, 16'hC516, 16'hBCD5, 16'hB4D4, 16'hAC53, 16'hBCD5, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hB515, 16'hB515, 16'hB4D5, 16'hB4D5, 16'hB515, 16'h730C, 16'h9410, 16'h83CF, 16'hA515, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hB557, 16'h9493, 16'h7B8F, 16'h9452, 16'h83CF, 16'hB597, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD16, 16'hAD16, 16'hAD57, 16'hAD57, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hB598, 16'hA4D5, 16'h9D15, 16'hAD97, 16'h6B4D, 16'h3104, 16'hC5D6, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9C0F, 16'hB491, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h9492, 16'h9492, 16'h9CD3, 16'hF79E, 16'hFFDF, 16'hCE59, 16'h7BCF, 16'h9492, 16'h9492, 16'h9492, 16'h9492,
        16'h9492, 16'h9492, 16'hA514, 16'hFFDF, 16'hD69A, 16'h8410, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h8C51, 16'h8C51, 16'hEF5D, 16'hEF5D, 16'h8410, 16'h9492, 16'h9492, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h8C51, 16'h9492, 16'h8C51, 16'h9492, 16'h9492, 16'h8410, 16'hAD55, 16'hA514, 16'hAD55, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65A, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hBCD3, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD5D7, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hC4D3, 16'hAC10, 16'hCD15, 16'hAC11, 16'hB451, 16'hC515, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC516, 16'hCD56, 16'hAC11, 16'hA451, 16'h9410, 16'hA4D4, 16'hAD56, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD15, 16'hAD15, 16'hAD16, 16'hAD15, 16'hAD16, 16'hACD4, 16'h834D, 16'h5800, 16'hB492, 16'hFF5D,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'h940F, 16'h000, 16'h3104, 16'h4186, 16'h880, 16'h8C91, 16'hA514, 16'h9C93, 16'hBDD7, 16'h7B4D, 16'h9BCF, 16'hCD57, 16'hC516, 16'hC516, 16'hBCD5, 16'hAC93, 16'hA412, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hB515, 16'hBD15, 16'hB4D5, 16'hB4D5, 16'hB515, 16'hACD4, 16'h624A, 16'hACD4, 16'h7B4D, 16'hAD56, 16'hAD57, 16'hAD57, 16'hAD57, 16'hAD57, 16'hB597, 16'h734E, 16'h9C94, 16'h7B8F,
        16'h9493, 16'hB598, 16'hAD57, 16'hB557, 16'hB557, 16'hB557, 16'hAD16, 16'hAD57, 16'hB557, 16'hB557, 16'hB557, 16'hB597, 16'hB597, 16'hB557, 16'hB598, 16'hB598, 16'h9CD4, 16'hAD57, 16'h9CD4, 16'h2000, 16'h9491, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h8ACB, 16'hD596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h9492, 16'hEF5D, 16'hFFDF, 16'hD69A, 16'h8410, 16'h8C51, 16'h8410, 16'h9492, 16'h9CD3, 16'h9492, 16'h8410, 16'hC618, 16'hFFDF, 16'hCE59, 16'h8C51, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'h9CD3, 16'h9492, 16'h8C51, 16'hAD55, 16'hEF5D, 16'hD69A, 16'h9492, 16'h9492, 16'h8410, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h9CD3, 16'h8C51, 16'h8C51, 16'h8C51, 16'h9CD3, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE18, 16'hE6DA, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBC92, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE18, 16'hD618, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hBCD3, 16'h9B4E, 16'hCD15, 16'hB451, 16'hB451, 16'hC4D4, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hB493, 16'hA3D0, 16'hA411, 16'h9C93, 16'hB556, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD15, 16'hAD15, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD16, 16'hB556, 16'h838E, 16'h4800, 16'h8B0B, 16'hE659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hB4D3, 16'h4943, 16'h2800, 16'h6248, 16'h4985, 16'h28C3, 16'h2142, 16'h9D13, 16'hAD55, 16'h9C93, 16'hBD96, 16'h6289, 16'hA3D0, 16'hCD56, 16'hC516, 16'hC516, 16'hBD15, 16'hAC53, 16'hA452, 16'hC516, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hB4D5, 16'hB4D5, 16'hBD16, 16'h93D0, 16'h6ACB, 16'hACD4, 16'h7B4D, 16'hB557, 16'hAD57, 16'hAD57, 16'hAD57, 16'hB598, 16'hA515, 16'h6B4D, 16'hAD56, 16'h6B0B, 16'hA515, 16'hB598, 16'hB597, 16'hB557, 16'hB597, 16'hAD57, 16'hA516, 16'hB598, 16'hB557, 16'hB597, 16'hB597, 16'hB597, 16'hB597, 16'hB598, 16'hB598, 16'hB598, 16'h9CD4, 16'hAD57, 16'h6B4E, 16'h6289, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD96, 16'h6800, 16'hDE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hA514, 16'h9492, 16'h8410, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hD69A, 16'hDEDB, 16'hF79E, 16'hD69A, 16'h8410, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hD69A, 16'h8410, 16'h9492, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8410, 16'h9492, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h9CD3, 16'h8C51, 16'h8C51, 16'h8C51, 16'h9492, 16'h8C51, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hD69A, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65A, 16'hE65A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC515, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE659, 16'hDE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD5D7, 16'h8249, 16'hCD15, 16'hB452, 16'hB452, 16'hC4D4, 16'hCD15, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC4D5, 16'h9B8F, 16'hAC52, 16'h9451, 16'hB556, 16'hB516, 16'hAD56,
        16'hAD56, 16'hAD56, 16'hAD16, 16'hAD15, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD16, 16'hAD16, 16'hB557, 16'h9C52, 16'h5186, 16'h4800, 16'hB4D2, 16'hF75C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hCD95, 16'h7B0A, 16'h000, 16'h5A08, 16'h82CB, 16'h82CA, 16'h7B0B, 16'h3945, 16'h1902, 16'h9D13, 16'hAD14, 16'h9C93, 16'hB555, 16'h6207, 16'hB493, 16'hCD57, 16'hC516, 16'hC516, 16'hC516, 16'hA412, 16'hAC52, 16'hC516, 16'hBD15, 16'hBD15, 16'hBD16, 16'hBD15, 16'hB515, 16'hB515, 16'hB515, 16'hB4D5, 16'hB515, 16'hBD16, 16'h72CB,
        16'h9451, 16'hA4D3, 16'h7B8E, 16'hB598, 16'hAD57, 16'hB557, 16'hB557, 16'hB598, 16'h7B8F, 16'h9453, 16'hA4D5, 16'h734D, 16'hB597, 16'hB597, 16'hB597, 16'hB557, 16'hB598, 16'hA4D5, 16'hA516, 16'hB598, 16'hB597, 16'hB598, 16'hB598, 16'hB598, 16'hB598, 16'hB598, 16'hBDD8, 16'hAD57, 16'h9CD4, 16'h9CD3, 16'h000, 16'hB554, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h8B8D, 16'h92CB, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8410, 16'h8C51, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h9CD3, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h8C51, 16'hC618, 16'hF79E, 16'hDEDB, 16'h9492, 16'h9492, 16'h8410, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8410, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'h9492, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD597, 16'hD618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'hCDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h828A, 16'hC4D4, 16'hB492, 16'hB451, 16'hC514, 16'hC515, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'h9B8F, 16'hB493, 16'h9410, 16'hB556, 16'hB556, 16'hB556, 16'hB556, 16'hB556, 16'hAD16, 16'hAD15, 16'hAD56, 16'hAD56, 16'hAD56, 16'hAD56, 16'hAD56, 16'hAD57, 16'hB557, 16'hAD15, 16'h7B4E, 16'h3800, 16'h58C1, 16'hBD14, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD5D7, 16'h830C, 16'h2000, 16'h38C2, 16'h7289, 16'h9B8D, 16'h8B0B, 16'hB450, 16'h8B4D, 16'h3103, 16'h3144, 16'h9C92, 16'hACD4, 16'hA4D3, 16'hB514, 16'h61C7, 16'hBCD4, 16'hCD57, 16'hC516, 16'hBD16, 16'hBD15, 16'h9BD0, 16'hB493, 16'hC516, 16'hBD15, 16'hBD16, 16'hBD16, 16'hBD15, 16'hB515, 16'hB516, 16'hB515, 16'hB4D5, 16'hBD16, 16'hAC94, 16'h49C7, 16'hB515, 16'h9C92, 16'h8C11, 16'hBD98, 16'hB557, 16'hB557, 16'hB598, 16'hA515, 16'h734E, 16'hB598, 16'h8C52, 16'h8C10, 16'hBDD8, 16'hB597, 16'hB598, 16'hB598, 16'hBD98, 16'h9493, 16'hB597, 16'hB598, 16'hB598, 16'hB598, 16'hB598, 16'hB598, 16'hB597, 16'hBDD8, 16'hBDD9, 16'hA516, 16'h8411, 16'h5ACB, 16'h6248, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h8B0B, 16'hBC51, 16'hF75D,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8C51, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hBDD7, 16'h8410, 16'h9CD3, 16'h8C51, 16'h9492, 16'h8C51, 16'h9492, 16'h8C51, 16'h9CD3, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'hAD55, 16'h9CD3, 16'h9CD3, 16'hBDD7, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hDE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'hCD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE659, 16'hD5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9BCF, 16'hB452, 16'hC4D4, 16'hAC10, 16'hCD15, 16'hC4D4, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD56,
        16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hD556, 16'hA3D0, 16'hAC92, 16'h9C11, 16'hACD4, 16'hB557, 16'hB556, 16'hB556, 16'hB556, 16'hAD56, 16'hA4D5, 16'hAD56, 16'hB556, 16'hB556, 16'hB557, 16'hB557, 16'hB557, 16'hAD57, 16'hB557, 16'hB557, 16'hA4D4, 16'h7B4D, 16'h2000, 16'h7207, 16'hC555, 16'hF75C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD618, 16'h8B8D, 16'h000, 16'h3902, 16'h5A07, 16'h830B, 16'h9BCD, 16'h8B4C, 16'hA40F, 16'hB4D2, 16'h9C50, 16'h2800, 16'h4A07, 16'h9C93, 16'hA4D4, 16'hACD4, 16'hAC93, 16'h7249, 16'hCD56, 16'hC556, 16'hC516, 16'hBD16, 16'hBCD4, 16'h8B8F, 16'hBCD4,
        16'hBD16, 16'hBD16, 16'hBD16, 16'hBD16, 16'hBD16, 16'hBD15, 16'hBD15, 16'hB515, 16'hB4D5, 16'hBD56, 16'h838E, 16'h734D, 16'hC5D8, 16'h8C10, 16'h9452, 16'hBDD8, 16'hB598, 16'hB598, 16'hBDD8, 16'h7BCF, 16'hA515, 16'hBD98, 16'h7B8F, 16'h9CD4, 16'hBDD8, 16'hB598, 16'hB598, 16'hBDD8, 16'hA515, 16'h9CD4, 16'hBDD8, 16'hB598, 16'hB598, 16'hB598, 16'hBDD8, 16'hA516, 16'h9D15, 16'hBE19, 16'hBE19, 16'h94D3, 16'h5ACB, 16'h6A8A, 16'hA491, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA450, 16'hC4D3, 16'hD596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8410, 16'h9CD3, 16'h8C51, 16'hAD55, 16'hDEDB, 16'hEF5D, 16'hEF5D, 16'hCE59, 16'h9492, 16'h9492, 16'h8C51, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hA514, 16'h8410, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hF79E, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD5D7, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'hBCD3, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69B, 16'hD5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD14, 16'h9B8F, 16'hCD15, 16'hAC10, 16'hCD15, 16'hC4D4, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hD557, 16'hB452, 16'h9BD0, 16'hAC52, 16'h9C92, 16'hBD97, 16'hB556, 16'hB556, 16'hB556, 16'hB557, 16'hAD15, 16'hB516, 16'hB556, 16'hB556, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hBD97, 16'hACD4, 16'h6ACC, 16'h000, 16'h6185, 16'hBD14, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9D, 16'hD618, 16'h8BCE, 16'h1800, 16'h2800, 16'h72CA, 16'h7289, 16'h9B8D, 16'hA40F, 16'h934C, 16'hAC50, 16'hAC50, 16'hC596, 16'hB513, 16'h40C1, 16'h628A, 16'h9492, 16'h9C92, 16'hACD4, 16'h93CF, 16'h8B0D, 16'hCD57, 16'hC556, 16'hBD16, 16'hC516, 16'hAC52, 16'h8B4E, 16'hBD16, 16'hBD16, 16'hBD16, 16'hBD16, 16'hBD16, 16'hBD16, 16'hBD16, 16'hBD16, 16'hB515, 16'hB515, 16'hB4D4, 16'h6289, 16'hAD15, 16'hC5D8, 16'h7B4D, 16'hA4D4, 16'hBDD9, 16'hB598, 16'hBDD8, 16'hAD15, 16'h9CD3, 16'hBDD8, 16'hAD56, 16'h734D, 16'hB597, 16'hB5D8, 16'hB598, 16'hBD98, 16'hBD98, 16'h8411, 16'hB597, 16'hBDD8, 16'hBD98, 16'hBD98, 16'hBDD9, 16'hB598, 16'h8412, 16'hBDD8, 16'hC65A, 16'hB597, 16'h738E, 16'h734D, 16'hB514, 16'hCDD7, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'hAC92, 16'hDDD7, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8410, 16'h9492, 16'h8C51, 16'h8410, 16'h9492, 16'h8C51, 16'h8410, 16'h9492, 16'h9492, 16'h8410, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hC618, 16'h9CD3, 16'h8C51, 16'h8C51, 16'hB596, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE18, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hBCD3, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hCD96, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hD5D7, 16'h828B, 16'hCD55, 16'hAC10, 16'hCD55, 16'hC4D4, 16'hCD56, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD57, 16'hC4D5, 16'h938F, 16'hB493, 16'h9C11, 16'hBD97, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hAD16, 16'hAD15, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hBD98, 16'hBD98, 16'hA4D4, 16'h7B4D, 16'h000, 16'h5942, 16'hA451, 16'hDE59, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5D, 16'hC595, 16'h834C, 16'h000, 16'h000, 16'h6A88, 16'h7ACA, 16'h7288, 16'h934C, 16'hB450, 16'h9B8D, 16'hAC10, 16'hAC51, 16'hBD14, 16'hD5D7, 16'hAC92, 16'h38C1, 16'h734C,
        16'h7B8E, 16'h9410, 16'hACD3, 16'h7ACB, 16'hAC11, 16'hCD57, 16'hC516, 16'hC516, 16'hC556, 16'h938F, 16'h9BD0, 16'hC556, 16'hBD16, 16'hBD16, 16'hBD16, 16'hBD16, 16'hBD16, 16'hBD16, 16'hBD16, 16'hB515, 16'hBD56, 16'h93D0, 16'h6B0C, 16'hC5D8, 16'hB556, 16'h6B0B, 16'hB597, 16'hBDD9, 16'hBDD9, 16'hB557, 16'h9493, 16'hB598, 16'hBDD9, 16'h9493, 16'h8C11, 16'hBDD9, 16'hBDD8, 16'hB598, 16'hBE19, 16'h9CD4, 16'h9493, 16'hC619, 16'hBDD8, 16'hBDD8, 16'hBDD9, 16'hC619, 16'h9493, 16'hA515, 16'hC65A, 16'hC619, 16'h8C11, 16'h6B0C, 16'hAD14, 16'hC596, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA410, 16'hE69A, 16'hBCD3, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8410, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h8410, 16'h9492, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hF79E, 16'hEF5D, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hE659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD96, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'hC555, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE659, 16'h7A49, 16'hC514, 16'hAC10, 16'hCD15, 16'hCD15, 16'hCD15, 16'hD556, 16'hD556, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hD556, 16'h9B4E, 16'hB493, 16'h9C10, 16'hB556, 16'hBD57, 16'hBD57, 16'hB557, 16'hB557, 16'hB556, 16'h9C93, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hB556, 16'hB597, 16'hB598, 16'hBD98, 16'hC5D8, 16'hAD15,
        16'h7B8F, 16'h3040, 16'h000, 16'h834B, 16'hC595, 16'hEF1B, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1B, 16'hBD54, 16'h728A, 16'h000, 16'h000, 16'h5A07, 16'h8B0B, 16'h82CA, 16'h9B8D, 16'h9B8D, 16'hA3CE, 16'h9B8D, 16'hAC50, 16'hB491, 16'hBD14, 16'hCDD7, 16'hCDD7, 16'hAC92, 16'h2800, 16'h7B4D, 16'h734D, 16'h838E, 16'h9C51, 16'h6A89, 16'hBCD4, 16'hCD57, 16'hC556, 16'hC556, 16'hBD15, 16'h624A, 16'hA452, 16'hC556, 16'hBD16, 16'hBD16, 16'hBD16, 16'hBD16, 16'hBD16, 16'hB4D4, 16'hBD16, 16'hBD16, 16'hBD15, 16'h628A, 16'h9C93, 16'hC5D8, 16'hA4D4, 16'h738E, 16'hBDD9, 16'hBDD9, 16'hBDD8, 16'h8C11, 16'hAD56, 16'hBDD9, 16'hBDD8, 16'h7B8E, 16'hAD16, 16'hBDD9, 16'hBDD8, 16'hBDD9, 16'hB597, 16'h7BD0, 16'hBDD8, 16'hBDD9, 16'hBDD9, 16'hBDD9,
        16'hC619, 16'hA515, 16'h8C52, 16'hC619, 16'hBDD8, 16'h8C51, 16'h8C10, 16'h9C51, 16'hF75D, 16'hD618, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC596, 16'hBD55, 16'hE659, 16'hBCD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hBDD7, 16'h9CD3, 16'h9492, 16'h9CD3, 16'hA514, 16'hC618, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hD5D7,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69B, 16'hC555, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hCD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'h8ACB, 16'hBC92, 16'hBC92, 16'hC4D4, 16'hCD55, 16'hC515, 16'hD556, 16'hCD56, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hCD56, 16'hD597, 16'hA3D0, 16'hA411, 16'hAC52, 16'hAC93, 16'hBD98, 16'hBD57, 16'hB557, 16'hB557, 16'hB557, 16'h9452, 16'hAD16, 16'hBD57, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hAD16, 16'hB557, 16'hBD98, 16'hB598, 16'hB598, 16'hBDD9, 16'hBDD9, 16'hB557, 16'h9492, 16'h5249, 16'h000, 16'h3800, 16'h938E, 16'hCDD6, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hE69A, 16'hA450, 16'h4942, 16'h000, 16'h3102, 16'h5A07, 16'h830A, 16'h934B, 16'h8B0B, 16'h934D,
        16'h934C, 16'h9B8D, 16'h9B8D, 16'hA3CF, 16'hB492, 16'hBD14, 16'hCDD7, 16'hCD96, 16'hCDD7, 16'hBD14, 16'h4944, 16'h628A, 16'h6ACA, 16'h5208, 16'h72CB, 16'h7ACB, 16'hCD56, 16'hC556, 16'hC556, 16'hCD57, 16'hA452, 16'h4184, 16'hACD3, 16'hC556, 16'hBD16, 16'hBD16, 16'hBD16, 16'hBD56, 16'hB4D4, 16'h834E, 16'hBD16, 16'hC557, 16'h93D0, 16'h62CC, 16'hBD97, 16'hC598, 16'h9452, 16'h8C51, 16'hC619, 16'hBDD8, 16'h83D0, 16'h9452, 16'hC5D9, 16'hBDD9, 16'hA4D5, 16'h7BCF, 16'hC5D9, 16'hBDD9, 16'hC619, 16'hC619, 16'h7BD0, 16'hAD56, 16'hC65A, 16'hBE19, 16'hBE19, 16'hC619, 16'hBDD8, 16'h8411, 16'hBDD8, 16'hBDD8, 16'h7BCF, 16'hB555, 16'h9C51, 16'hDE9A, 16'hF75D, 16'hCDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h8B4C, 16'hF6DC, 16'hBC92, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hF79E, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD5D7, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hBD13, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC514, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hB450, 16'hB451, 16'hBC92, 16'hCD15, 16'hD556, 16'hC4D4, 16'hCD56, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD597, 16'hB453, 16'hA3D0, 16'hB4D4, 16'h9411, 16'hBD98, 16'hBD57, 16'hB597, 16'hB557, 16'hBD97, 16'h9C52, 16'hA4D4, 16'hBD98, 16'hB557,
        16'hB597, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hB557, 16'hAD15, 16'hB598, 16'hB598, 16'hB598, 16'hBD98, 16'hBD98, 16'hBDD9, 16'hC5D9, 16'hBD98, 16'hAD15, 16'h83D0, 16'h49C8, 16'h000, 16'h48C0, 16'h93CF, 16'hC596, 16'hEF1B, 16'hFFDE, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1B, 16'hC595, 16'h7B0B, 16'h40C0, 16'h000, 16'h2903, 16'h6248, 16'h6A88, 16'h7AC9, 16'h8B4B, 16'h934C, 16'h938C, 16'h9B8D, 16'hA3CE, 16'hA3CE, 16'h938E, 16'hC514, 16'hBD13, 16'hCDD7, 16'hCDD6, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'h838D, 16'h4145, 16'h6249, 16'h6289, 16'h4102, 16'h9BCF, 16'hCD57, 16'hC556, 16'hC556, 16'hC516, 16'h6ACB, 16'h7B4D, 16'hBD15, 16'hC516, 16'hBD16, 16'hBD16, 16'hBD16, 16'hC557, 16'h9C11, 16'h834D, 16'hC557, 16'hBD56, 16'h628A, 16'h9C93, 16'hC5D8, 16'hB556, 16'h6B0C, 16'hB597, 16'hC619, 16'h7B8F, 16'h7BD0, 16'hC619, 16'hBDD9, 16'hBDD8,
        16'h7B8E, 16'hA4D5, 16'hC619, 16'hC5D9, 16'hBE19, 16'h7BCF, 16'h9493, 16'hCE5A, 16'hC61A, 16'hBE19, 16'hC61A, 16'hCE5A, 16'h83D0, 16'hA514, 16'hAD56, 16'h83CF, 16'hD618, 16'hBD14, 16'hC596, 16'hFFDF, 16'hCE18, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h8B4B, 16'hDE59, 16'hDE59, 16'hBCD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hD5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCDD7, 16'hDE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD96, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hBCD3, 16'hB493, 16'h8B0B, 16'hCD15, 16'hD597, 16'hC4D4, 16'hCD15, 16'hD556, 16'hD556, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hD556, 16'hD557, 16'hCD15, 16'h934E, 16'hBCD5, 16'h93D0, 16'hBD57, 16'hBD98, 16'hBD98, 16'hBD97, 16'hBD97, 16'hAD15, 16'h8C11, 16'hBD57, 16'hBD97, 16'hBD97, 16'hBD57, 16'hBD57, 16'hBD57, 16'hBD57, 16'hB557, 16'hBD98, 16'hAD16, 16'hAD15, 16'hBDD8, 16'hBDD8, 16'hBD98, 16'hBD98, 16'hBDD8, 16'hBDD8, 16'hBDD9, 16'hC5D9, 16'hC5D9, 16'hBD98, 16'hA515, 16'h83D0, 16'h49C7, 16'h000, 16'h4040, 16'h834C, 16'hCDD7, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79D, 16'hDE99, 16'hA4D1, 16'h51C5,
        16'h000, 16'h2840, 16'h49C6, 16'h51C6, 16'h7289, 16'h7288, 16'h72C9, 16'h830B, 16'h8B4C, 16'h8B4C, 16'h938D, 16'h9B8D, 16'hAC50, 16'h9BCE, 16'hBCD3, 16'hB4D3, 16'hCDD7, 16'hCDD7, 16'hCDD6, 16'hCDD7, 16'hCDD7, 16'hD618, 16'h9C10, 16'h4103, 16'h730B, 16'h834C, 16'h4903, 16'hB493, 16'hCD57, 16'hC556, 16'hCD57, 16'hAC92, 16'h4144, 16'h8B8E, 16'hC516, 16'hC516, 16'hC556, 16'hC556, 16'hBD56, 16'hC556, 16'h72CC, 16'h9C11, 16'hCD98, 16'hAC93, 16'h730D, 16'hBD97, 16'hC5D8, 16'h9C93, 16'h8411, 16'hBDD8, 16'h734F, 16'h8411, 16'hBDD9, 16'hC619, 16'hC61A, 16'hA514, 16'h734E, 16'hC5D9, 16'hCE5A, 16'hBDD8, 16'h738E, 16'h9452, 16'hCE9B, 16'hCE9B, 16'hCE5A, 16'hC61A, 16'hC619, 16'h8410, 16'h8C10, 16'hA492, 16'hBD14, 16'hE69A, 16'hBD55, 16'hBD55, 16'hFFDF, 16'hF75D, 16'hC596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hA40F, 16'hC596, 16'hFFDF, 16'hB4D2, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD5D7, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hEF1D, 16'hB492, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hDE18, 16'hE659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC514, 16'hDE18, 16'h934D, 16'hBC92, 16'hDD97, 16'hCD15, 16'hBC52, 16'hD556, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hD556, 16'hD557,
        16'h9B8F, 16'hB453, 16'hA411, 16'hACD4, 16'hC5D8, 16'hBD98, 16'hBD98, 16'hC5D8, 16'hB556, 16'h9452, 16'hA493, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD97, 16'hBD97, 16'hBD97, 16'hBD97, 16'hBD98, 16'h9492, 16'hA4D4, 16'hBDD8, 16'hBDD9, 16'hBDD9, 16'hBDD9, 16'hBDD9, 16'hBDD9, 16'hC5D9, 16'hC5D9, 16'hC5D9, 16'hC61A, 16'hC5D9, 16'hBDD8, 16'hAD56, 16'h8C10, 16'h5209, 16'h1800, 16'h3800, 16'h940F, 16'hCE17, 16'hEF1C, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79D, 16'hDE99, 16'hB513, 16'h72CA, 16'h2800, 16'h000, 16'h3104, 16'h6248, 16'h5A07, 16'h5A06, 16'h6A48, 16'h7AC9, 16'h834C, 16'h7ACA, 16'h8B4C, 16'h938D, 16'h938D, 16'hAC50, 16'hB491, 16'h8B0C, 16'hC513, 16'hB4D2, 16'hC596, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hCDD6, 16'hB514, 16'h6248, 16'h4984, 16'h93CF, 16'h8B4D, 16'h6A8A, 16'hCD56, 16'hC556, 16'hC556, 16'hCD56, 16'h8B8E, 16'h7B4C, 16'h8BCE, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC557, 16'hB4D4, 16'h59C8, 16'hB4D5, 16'hCD97, 16'h7B4D,
        16'h9452, 16'hC5D8, 16'hBD56, 16'h734D, 16'hAD15, 16'h8C11, 16'h8410, 16'hBDD8, 16'hC5D9, 16'hB556, 16'hB556, 16'h734D, 16'hAD56, 16'hCE5A, 16'hA4D4, 16'h7B8D, 16'hA514, 16'hD69B, 16'hCE5A, 16'hB597, 16'hAD16, 16'h9CD4, 16'h5A8B, 16'h8BCF, 16'hDE9A, 16'hEF1D, 16'hEF1C, 16'hAD13, 16'hB514, 16'hFFDF, 16'hFFDF, 16'hD5D7, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hA410, 16'hB4D2, 16'hFFDF, 16'hCD97, 16'hC555, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hCD55, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hC555, 16'hD618, 16'hFFDF, 16'hFFDF, 16'hE659, 16'hDDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCDD7, 16'hE659, 16'hB4D3, 16'hA38F, 16'hDD97, 16'hD556, 16'hBC52, 16'hC4D4, 16'hD597, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hD597, 16'hB452, 16'h9B8F, 16'hC515, 16'h93D0, 16'hC598, 16'hC5D8, 16'hC5D8, 16'hC5D8, 16'hBD97, 16'hB515, 16'hA493, 16'hAD15, 16'hC5D9, 16'hC598, 16'hC5D8, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD98, 16'hC5D8, 16'hB556, 16'h8C51, 16'hAD16, 16'hAD56, 16'hBD98, 16'hC5D9, 16'hC5D9, 16'hBDD9, 16'hC5D9, 16'hC5D9, 16'hC5D9, 16'hC619, 16'hBD98, 16'hBD98, 16'hD65B, 16'hDE9B, 16'hCE19, 16'hAD15, 16'h8C10, 16'h2000, 16'h1000, 16'h59C4, 16'h9C0E, 16'hC595,
        16'hDE58, 16'hDE59, 16'hD618, 16'hBD54, 16'h9C4F, 16'h6AC9, 16'h3900, 16'h000, 16'h1000, 16'h3985, 16'h5207, 16'h6247, 16'h5206, 16'h6247, 16'h6A88, 16'h938C, 16'h8B4B, 16'h7B0A, 16'h834B, 16'h938D, 16'h938D, 16'hA40F, 16'hBC91, 16'h8B4C, 16'hBCD2, 16'hB491, 16'hC555, 16'hCDD7, 16'hCDD7, 16'hC596, 16'hBD54, 16'hA410, 16'h6A48, 16'h4985, 16'h8B8E, 16'hBD54, 16'hBD54, 16'h5184, 16'h9C11, 16'hCD97, 16'hC556, 16'hCD57, 16'hAC92, 16'h6A89, 16'hA451, 16'h8B8E, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hCD57, 16'h93CF, 16'h6A8B, 16'hC557, 16'hB515, 16'h628A, 16'hB556, 16'hC5D8, 16'h8BD0, 16'h734D, 16'hC5D7, 16'hA4D3, 16'hAD14, 16'h9410, 16'hACD3, 16'hA4D3, 16'h7B8E, 16'h8C10, 16'hC5D7, 16'hBD55, 16'h9451, 16'hC5D7, 16'hC5D7, 16'h9C92, 16'h8C10, 16'h8C10, 16'hA492, 16'h93CF, 16'hAD13, 16'hFF9E, 16'hFFDF, 16'hD659, 16'h940F, 16'hCDD7, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'hC554, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hA410, 16'hBCD3, 16'hFFDF, 16'hEF1C, 16'hAC10, 16'hFF9E,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hA514, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hD596, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hBCD2, 16'hE69A, 16'hFFDF, 16'hEF1B, 16'hC515, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'hC555, 16'hE69A, 16'h930C, 16'hDD97,
        16'hDD57, 16'hCD14, 16'hA3CF, 16'hD556, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hD516, 16'h8ACC, 16'hCD15, 16'hA451, 16'hB515, 16'hCE19, 16'hC5D9, 16'hC5D8, 16'hC5D8, 16'hACD4, 16'hCE19, 16'h9C52, 16'hC598, 16'hC5D9, 16'hC5D8, 16'hC5D8, 16'hC598, 16'hBD98, 16'hBD98, 16'hBD98, 16'hC5D9, 16'hA4D4, 16'h8C10, 16'hB557, 16'h9C93, 16'hA515, 16'hBD98, 16'hC61A, 16'hCE1A, 16'hCE1A, 16'hCE1A, 16'hCE1A, 16'hCE1A, 16'hB556, 16'hA4D4, 16'hC5D9, 16'hD65B, 16'hDE9C, 16'hDE9C, 16'hC5D9, 16'hA515, 16'h7BCE, 16'h730B, 16'h51C5, 16'h3880, 16'h3000, 16'h38C0, 16'h000, 16'h800, 16'h1800, 16'h3144, 16'h49C6, 16'h5206, 16'h5A07, 16'h72C9, 16'h6A47, 16'h6A88, 16'h5A06, 16'h8B8C, 16'h834B, 16'h7B0A, 16'h8B4C, 16'hA40E, 16'h9BCE, 16'hAC0F, 16'hAC50, 16'h938D, 16'hAC50, 16'hBCD3, 16'hC554, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hC5D6, 16'hACD2, 16'hA451, 16'hAC92, 16'hBD55, 16'hD618, 16'hDE59, 16'hA451, 16'h6207, 16'hC515, 16'hC556, 16'hC557, 16'hC515, 16'h5A48, 16'h5A08,
        16'h6A89, 16'h9C10, 16'hCD57, 16'hC556, 16'hC556, 16'hC557, 16'hBD15, 16'h59C7, 16'h93D0, 16'hCDD8, 16'h8BD0, 16'h734D, 16'hC5D8, 16'hACD4, 16'h49C7, 16'hBD55, 16'hFFDF, 16'hFF9F, 16'hF75E, 16'hF75E, 16'hEF1C, 16'h83CF, 16'h9450, 16'hF79D, 16'hF79E, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hDE9A, 16'hDE9A, 16'hEF1C, 16'hF75D, 16'hD618, 16'hCD96, 16'hFF9E, 16'hEEDB, 16'hAC92, 16'hA451, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD95, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'h934D, 16'hCDD7, 16'hFFDF, 16'hFF9F, 16'hAC10, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'hBDD7, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8410, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hDE18, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hAC10, 16'hF71C, 16'hFFDF, 16'hC514, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hBCD3, 16'hFF5D, 16'hA3CF, 16'hBC93, 16'hDD97, 16'hDD57, 16'hABCF, 16'hC4D3, 16'hDD97, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hDD97, 16'hABD0, 16'hAC11, 16'hCD16, 16'h9C10, 16'hD619, 16'hCDD9, 16'hCDD9, 16'hCE19, 16'hAD15, 16'hCE18, 16'hDE9A, 16'h8BD0, 16'hC598, 16'hC5D9, 16'hC598, 16'hC5D8, 16'hC5D8, 16'hC598, 16'hC5D8, 16'hC5D9, 16'hC5D8, 16'h9452, 16'hA515, 16'hC5D9, 16'hAD15, 16'h8C51, 16'h9493, 16'hAD55, 16'hC5D8, 16'hCE19, 16'hCE19,
        16'hCE1A, 16'hD65A, 16'hB556, 16'h7B8F, 16'hA4D4, 16'hC5D8, 16'hDE9B, 16'hCE5A, 16'hC618, 16'hDE9A, 16'hBD54, 16'h4140, 16'h83CE, 16'hA4D2, 16'h7B4C, 16'h3984, 16'h4A06, 16'h41C5, 16'h4185, 16'h5A07, 16'h51C6, 16'h6248, 16'h6288, 16'h7B0A, 16'h6247, 16'h6A88, 16'h7B0B, 16'h7B0B, 16'h938D, 16'hA40F, 16'h9BCD, 16'hA40F, 16'hAC50, 16'hAC50, 16'hA410, 16'hC554, 16'hBD14, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCE17, 16'hD617, 16'hD618, 16'hCDD7, 16'hCDD7, 16'hC596, 16'h5185, 16'hAC92, 16'hCD97, 16'hC556, 16'hCD97, 16'h838D, 16'h6ACA, 16'hAC92, 16'h3902, 16'hA452, 16'hCD97, 16'hC556, 16'hC556, 16'hCD57, 16'h9C11, 16'h38C3, 16'hBD15, 16'hB514, 16'h5A48, 16'hAD15, 16'hB556, 16'h628B, 16'hBD96, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h9C91, 16'h9410, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD95, 16'hA410, 16'hD5D7, 16'hC596, 16'hBD14, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE19, 16'hC555, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hBD14, 16'hAC92, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hCD95, 16'hCD95, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h7BCF, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8C51, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hDE18, 16'hF75E, 16'hFFDF, 16'hE69B,
        16'hB411, 16'hF6DC, 16'hCD96, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD96, 16'hEE9B, 16'hE659, 16'h9B4D, 16'hE597, 16'hDD97, 16'hCCD4, 16'hA38E, 16'hDD97, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hD597, 16'hD557, 16'hDD97, 16'hCCD5, 16'h8249, 16'hCD15, 16'hAC11, 16'hBD15, 16'hD61A, 16'hCE19, 16'hCE19, 16'hC5D8, 16'hA4D3, 16'hF75E, 16'hD619, 16'h8BD0, 16'hC598, 16'hCDD9, 16'hC5D9, 16'hC5D9, 16'hC5D9, 16'hC5D9, 16'hC5D9, 16'hC5D9, 16'hC619, 16'h8C51, 16'hAD56, 16'hC5D8, 16'hE6DC, 16'hC5D8, 16'h9C93, 16'h9C92, 16'h9C92, 16'h9C92, 16'hBDD7, 16'hE71C, 16'hE71C, 16'hD65A, 16'hBDD7, 16'hB515, 16'h9C92, 16'hAD55, 16'hF75D, 16'hCE17, 16'h2800, 16'h9450, 16'hC5D6, 16'h9C50, 16'h730A, 16'h5A47, 16'h28C1, 16'h5206, 16'h6247, 16'h5A47, 16'h6A89, 16'h5A06, 16'h72CA, 16'h6A48, 16'h6248, 16'h7B0A, 16'h834C, 16'h834C, 16'hAC50, 16'h9BCD, 16'hAC4F, 16'hA40E, 16'hBCD1, 16'h93CE, 16'hC554, 16'hC595, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7,
        16'hCDD7, 16'hCDD7, 16'hD617, 16'h8BCE, 16'h7289, 16'hC555, 16'hC556, 16'hCD97, 16'hA451, 16'h3902, 16'hB514, 16'hAC93, 16'h5A07, 16'hC556, 16'hCD57, 16'hC556, 16'hCD57, 16'hBD15, 16'h4145, 16'h834E, 16'hC556, 16'h6ACA, 16'h8BD0, 16'hBD56, 16'h5A48, 16'h838D, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hC596, 16'h7B0B, 16'hAD13, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hFFDF, 16'hFF9F, 16'hF75D, 16'hCE18, 16'h940F, 16'hACD2, 16'hDE59, 16'hDE5A, 16'hEF1D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE5A, 16'hBCD3, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hD618, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE18, 16'hBD13, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8C51, 16'h9492, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h8C51, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hEE9A, 16'hEEDB, 16'hFFDF, 16'hEE9B, 16'hBC52, 16'hB410, 16'hD5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hCD96, 16'hFFDF, 16'hA3CF, 16'hC493, 16'hE5D8, 16'hE597, 16'hABD0, 16'hBC93, 16'hDD98, 16'hD557, 16'hD597, 16'hD557, 16'hD597, 16'hD597, 16'hD597, 16'hD557, 16'hDD97, 16'h9B8E, 16'h9B4E, 16'hDD97, 16'h9BCF, 16'hCE19, 16'hD65A, 16'hCE19, 16'hD65A, 16'hB555, 16'hCE18, 16'hFFDF, 16'hD659, 16'h9411, 16'hBD97, 16'hCE1A, 16'hCDD9, 16'hC5D9, 16'hC5D9,
        16'hC5D9, 16'hC5D9, 16'hCE1A, 16'hC5D8, 16'h8C51, 16'h9C93, 16'hEF5D, 16'hFFDF, 16'hFF9F, 16'hF75D, 16'hEF5D, 16'hF79E, 16'hFFDF, 16'hFF9F, 16'hEF1C, 16'hE6DC, 16'hE71C, 16'hCE59, 16'hC5D7, 16'hF75D, 16'hF79E, 16'h6B0B, 16'h6B0B, 16'hCDD7, 16'h9C91, 16'h72C9, 16'hA44F, 16'h940F, 16'h49C6, 16'h4985, 16'h6247, 16'h5A47, 16'h6247, 16'h6AC9, 16'h6A88, 16'h6247, 16'h8B4C, 16'h8B4C, 16'h834C, 16'hA44F, 16'h93CD, 16'h9BCE, 16'h9BCE, 16'hB491, 16'hA40F, 16'hC514, 16'hCD96, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hACD2, 16'h4902, 16'hB4D3, 16'hC556, 16'hCD97, 16'hBCD4, 16'h4984, 16'h940F, 16'hCDD7, 16'h8BCF, 16'h72CB, 16'hCD97, 16'hC556, 16'hC556, 16'hC556, 16'h7B4D, 16'h51C7, 16'hACD3, 16'h93CF, 16'h6ACB, 16'h9C51, 16'h51C6, 16'h9C91, 16'hE6DA, 16'hC596, 16'hB554, 16'hA491, 16'h8BCE, 16'h9C91, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'hC596, 16'hB4D3, 16'hACD2, 16'hACD2, 16'hE6DB, 16'hFF9E,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD617, 16'hBD14, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE659, 16'hBC92, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hB596, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hF71C, 16'hF71C, 16'hF71C, 16'hBC93, 16'hA38F, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hBCD3, 16'hFF5D, 16'hE6DB, 16'h9B4D, 16'hDD97, 16'hE5D8, 16'hD515, 16'hA38D, 16'hD556, 16'hDD98, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD98, 16'hD515, 16'h8249, 16'hAC11, 16'hBC92, 16'hBD14, 16'hDE5A, 16'hCE19, 16'hD65A, 16'hD619, 16'hA411, 16'hEF1C, 16'hFFDF, 16'hE6DB, 16'h9C92, 16'hA4D4, 16'hC5D9, 16'hD65A, 16'hD61A, 16'hCE1A, 16'hCE1A, 16'hCE1A, 16'hCE1A, 16'hCE19, 16'h8410, 16'hA4D3, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1D, 16'hCE18, 16'hC5D7, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hCE17, 16'h800, 16'hAD54, 16'hBD95, 16'h5A06, 16'hA450, 16'hB513, 16'hB513, 16'h6ACA, 16'h2880, 16'h5A07, 16'h5A47, 16'h6247, 16'h6248, 16'h6247, 16'h93CE, 16'h93CD, 16'h8B4C, 16'h9C0E, 16'h9C0F, 16'h9BCE, 16'hA40F, 16'hAC50, 16'hAC50,
        16'hBCD2, 16'hCD95, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCD96, 16'h6A48, 16'h834C, 16'hC556, 16'hCD56, 16'hB4D3, 16'h5184, 16'h8B8E, 16'hC5D7, 16'hC596, 16'h6A89, 16'h9C11, 16'hCD97, 16'hC556, 16'hCD97, 16'h838E, 16'h49C6, 16'h8BCF, 16'h730B, 16'h1000, 16'h5A47, 16'h62C9, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hE6DB, 16'hDEDB, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5C, 16'hE69A, 16'hD618, 16'hC555, 16'hD618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD5D7, 16'hC514, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hF79E, 16'h9CD3, 16'h8410, 16'h8410, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hB492, 16'hA38E, 16'hEE9A, 16'hF71C, 16'hFF9E, 16'hFFDF, 16'hE659, 16'hDE18, 16'hFFDF, 16'hBCD3, 16'hC493, 16'hE5D8, 16'hDD98, 16'hCCD3, 16'hB3D0, 16'hDD97, 16'hDD98, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD98, 16'hDD98, 16'hD598, 16'hE598, 16'hBC12, 16'h6946, 16'h9B4E, 16'hB411, 16'hCD97,
        16'hDE9B, 16'hD65A, 16'hD65A, 16'hCD97, 16'hB514, 16'hFF9F, 16'hFFDF, 16'hF79E, 16'hBD96, 16'h9C51, 16'hACD4, 16'hC5D8, 16'hD65A, 16'hD65B, 16'hD65B, 16'hCE5B, 16'hCE5B, 16'hCE5A, 16'hAD15, 16'h9CD2, 16'hC618, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h6288, 16'h734C, 16'hCE18, 16'hA4D3, 16'h6248, 16'hAC91, 16'hB512, 16'hB4D2, 16'h838C, 16'h1000, 16'h5206, 16'h6248, 16'h72C9, 16'h72C9, 16'h8B4C, 16'hA44F, 16'h834B, 16'h938D, 16'hAC90, 16'h938D, 16'hB491, 16'hB491, 16'hBCD2, 16'hC514, 16'hCD96, 16'hCDD6, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'h938E, 16'h4903, 16'hC555, 16'hCDD7, 16'hA451, 16'h4080, 16'h9410, 16'hC5D7, 16'hCE18, 16'hA451, 16'h6A89, 16'hC515, 16'hC557, 16'hCD96, 16'h93D0, 16'h1000, 16'h6289, 16'h6289, 16'h734C, 16'hA4D2, 16'hCE17, 16'hF79D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hEF5C, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hEF1C, 16'hDE18, 16'hDDD8, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h9492, 16'h8C51, 16'hDEDB, 16'hFFDF, 16'hC618, 16'h8410,
        16'h9CD3, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h8C51, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hA3CE, 16'hDD97, 16'hDDD7, 16'hCD14, 16'hD5D7, 16'hDDD7, 16'hB3D0, 16'hF71D, 16'hF6DC, 16'h9B0C, 16'hDD56, 16'hE5D9, 16'hE598, 16'hC493, 16'hBC51, 16'hE598, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD56, 16'h9B0C, 16'hAB8E, 16'hAB8F, 16'h9B4E, 16'hD597, 16'hE69B, 16'hDE9A, 16'hDE9B, 16'hC556, 16'hB4D4, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hCE18, 16'hA4D3, 16'h9452, 16'hA4D4, 16'hB596, 16'hC619, 16'hCE19, 16'hC619, 16'hCE1A, 16'hC5D9, 16'hA514, 16'hAD14, 16'hAD14, 16'hB555, 16'hC5D7, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD96, 16'h000, 16'hB554, 16'hCE18, 16'hB554, 16'h49C5, 16'hA490, 16'h9C4F, 16'hA44F, 16'h8B8D, 16'h1800, 16'h4184, 16'h72C9,
        16'h834B, 16'h834B, 16'hA44F, 16'h8B8C, 16'h93CD, 16'hB4D1, 16'h8B8D, 16'hBCD2, 16'hB491, 16'hCD95, 16'hCD95, 16'hD5D6, 16'hCDD7, 16'hCDD7, 16'hCDD6, 16'hCDD6, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'h9BCF, 16'h50C1, 16'hBD14, 16'hC595, 16'h72CA, 16'h6249, 16'hACD3, 16'hC5D7, 16'hCE18, 16'hB514, 16'h51C6, 16'hAC52, 16'hCD57, 16'hCD56, 16'h93CF, 16'h2800, 16'h834D, 16'h49C6, 16'h62C9, 16'hA4D2, 16'hBD95, 16'hBD95, 16'hC5D7, 16'hBD96, 16'hC5D7, 16'hB554, 16'hA4D2, 16'hA4D3, 16'hB554, 16'hBDD7, 16'hD659, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hF75D, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hCE59, 16'hB596, 16'hB596, 16'hC618, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8C51, 16'h8410, 16'hD69A, 16'hEF5D, 16'h8410, 16'h9492, 16'h8410, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8C51, 16'h8C51, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hAC0F, 16'hF71C, 16'hFF5D, 16'hE69A, 16'hE659, 16'hCD14, 16'hBC91, 16'hE618, 16'hCCD4, 16'h9A8B, 16'hE597, 16'hE5D8, 16'hE598, 16'hC492, 16'hBC11,
        16'hDD97, 16'hE5D8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hE5D8, 16'hC493, 16'hA34D, 16'hC452, 16'hB411, 16'h9B4E, 16'hBC93, 16'hCD97, 16'hDE5A, 16'hE69A, 16'hCD96, 16'hC556, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71B, 16'hC5D7, 16'hB514, 16'h9C92, 16'h9410, 16'h9C91, 16'h9450, 16'h9C92, 16'hAD14, 16'hA4D2, 16'hB555, 16'hD69A, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h5206, 16'h7B4C, 16'hC5D7, 16'hC5D7, 16'hC5D6, 16'h6ACA, 16'h8BCD, 16'hA450, 16'h9C0F, 16'h940E, 16'h51C6, 16'h3902, 16'h8B8C, 16'h93CD, 16'h9C0E, 16'h9C0E, 16'h938D, 16'hBCD2, 16'hA450, 16'hAC91, 16'hD5D6, 16'hCD96, 16'hD5D7, 16'hCDD7, 16'hCDD6, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hAC91, 16'h5144, 16'h9C0F, 16'h9C50, 16'h4982, 16'h834D, 16'hBD96, 16'hC5D8, 16'hCE18, 16'hBD55, 16'h6289, 16'h8B8E, 16'hC515, 16'hBD15, 16'h834D, 16'h4943, 16'h9451, 16'hC5D7, 16'h9450, 16'h49C5, 16'h838D,
        16'h8B8E, 16'h7B0C, 16'h72CB, 16'h5A48, 16'h5207, 16'h838D, 16'h9C10, 16'h8BCF, 16'h9410, 16'h8BCF, 16'h6ACB, 16'h7B4D, 16'hAD14, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h9CD3, 16'h8410, 16'h8C51,
        16'h8C51, 16'h8C51, 16'h8410, 16'hC618, 16'hFFDF, 16'hCE59, 16'h8410, 16'h9492, 16'hAD55, 16'h9CD3, 16'h8C51, 16'h8C51, 16'h9CD3, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8C51, 16'h8C51, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD5D7, 16'hABCF, 16'hE659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE619, 16'hE619, 16'hF6DC, 16'hC4D3, 16'h9209, 16'hD515, 16'hE5D8, 16'hEDD9, 16'hC493, 16'hBC10, 16'hDD97, 16'hE5D8, 16'hDD98, 16'hE598, 16'hE5D8, 16'hE598, 16'hE598, 16'hEDD8, 16'hAB8E, 16'hC493, 16'hEDD8, 16'hBC93, 16'hB451, 16'hBC93, 16'hB4D3, 16'hBD15, 16'hC515, 16'hC514, 16'hB492, 16'hD5D7, 16'hF71C, 16'hFF9E, 16'hFFDE, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hEF5D, 16'hF75D, 16'hF75D, 16'hE71C, 16'hF75D, 16'hF79D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB555, 16'h000,
        16'hB555, 16'hC617, 16'hC5D7, 16'hCE17, 16'h8BCE, 16'h6A89, 16'hAC90, 16'h8BCD, 16'h9C0F, 16'h7B0A, 16'h2800, 16'hA44F, 16'hBD13, 16'hAC50, 16'hAC90, 16'hA450, 16'hBD13, 16'h9C0F, 16'hD5D6, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'h9C0F, 16'h2800, 16'h59C5, 16'h6A89, 16'h7B4C, 16'hACD3, 16'hC5D7, 16'hC5D8, 16'hCE18, 16'hB555, 16'h72CA, 16'h8B8D, 16'hA451, 16'h93CF, 16'h5207, 16'h6ACB, 16'hAD14, 16'hC5D7, 16'hC618, 16'hAD54, 16'h5A48, 16'hACD3, 16'hC556, 16'hBD15, 16'hC556, 16'hBD55, 16'h7B4D, 16'hA492, 16'hC597, 16'hBD56, 16'hACD3, 16'h9C51, 16'h838E, 16'h6ACB, 16'h7B4D, 16'h6289, 16'hAD13, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hD69A, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h8C51, 16'h9492, 16'h8C51, 16'h8410, 16'h9492, 16'h9492, 16'h8C51, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8C51, 16'h9492, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hB3CF,
        16'hBC51, 16'hDE18, 16'hF71C, 16'hEE9B, 16'hDD96, 16'hFF5E, 16'hFF9E, 16'hDDD7, 16'hA30C, 16'hAB4E, 16'hD515, 16'hE598, 16'hC452, 16'hB3D0, 16'hDD57, 16'hE5D9, 16'hE5D8, 16'hE598, 16'hE598, 16'hE598, 16'hEDD9, 16'hDD56, 16'h930D, 16'hD556, 16'hF69A, 16'hCD55, 16'hC4D4, 16'hCD56, 16'hE65A, 16'hDE19, 16'hDE19, 16'hE69B, 16'hEEDC, 16'hE69A, 16'hE69A, 16'hEEDB, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71B, 16'h4983, 16'h83CE, 16'hCE18, 16'hC5D7, 16'hC5D7, 16'hCE18, 16'hA4D2, 16'h5A06, 16'hAC91, 16'h93CE, 16'h838C, 16'h8B8C, 16'h000, 16'hA450, 16'hD617, 16'hC595, 16'hC554, 16'hC555, 16'hC554, 16'hC555, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD6, 16'hCDD6, 16'hD617, 16'hC555, 16'h6ACA, 16'h000, 16'h7B4C, 16'hA492, 16'hB555, 16'hCE18, 16'hCE18, 16'hC5D7, 16'hC596, 16'hACD3, 16'h5207,
        16'h7289, 16'h7ACB, 16'h5A08, 16'h6B0B, 16'hA4D3, 16'hC5D7, 16'hC5D8, 16'hBDD7, 16'hC5D7, 16'hC5D7, 16'h8C0F, 16'h5206, 16'hB514, 16'hBD55, 16'hB514, 16'hBD55, 16'hB514, 16'hBD56, 16'hB514, 16'h7B0C, 16'h62CB, 16'h9C52, 16'hA493, 16'h9C52, 16'h9C52, 16'hA4D4, 16'h5A48, 16'hA4D2, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8C51, 16'h8410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'h9CD3, 16'h738E, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h8410, 16'h9492, 16'h8C51, 16'hC618, 16'hD69A, 16'hAD55, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'hA514, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h7BCF, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hDE59, 16'hBC92, 16'hBC91, 16'hD554, 16'hD514, 16'hCCD2, 16'hDDD7, 16'hEE9A, 16'hDDD7, 16'hCCD4, 16'hB38F, 16'hA2CC, 16'hBB8F, 16'hB34E, 16'h9A4A, 16'hC493, 16'hE598, 16'hEDD9, 16'hEDD9, 16'hEDD9, 16'hE5D8, 16'hEDD9, 16'hD515, 16'h9B0C, 16'hCD15, 16'hF69B, 16'hDDD8, 16'hB452, 16'hCCD4, 16'hEE9B, 16'hEEDB, 16'hF71C, 16'hF71D, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C,
        16'hE6DB, 16'hD659, 16'hB595, 16'h9C92, 16'hAD14, 16'hC5D6, 16'hBD95, 16'hC5D7, 16'hDE9A, 16'h8BCE, 16'h2840, 16'hB595, 16'hC618, 16'hC5D7, 16'hC5D7, 16'hCE18, 16'hBD95, 16'h4985, 16'h72CA, 16'h834C, 16'hA450, 16'h93CD, 16'h1800, 16'hA491, 16'hD617, 16'hCDD6, 16'hCDD6, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD6, 16'hCDD7, 16'hD5D7, 16'hB4D3, 16'h5984, 16'h728A, 16'hC555, 16'hDE59, 16'hE65A, 16'hD659, 16'hCE18, 16'hCE18, 16'hB555, 16'h838E, 16'h5A48, 16'h834D, 16'h9410, 16'h9C92, 16'hB555, 16'hC5D7, 16'hC618, 16'hC5D7, 16'hBDD7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hAD13, 16'h3943, 16'h6289, 16'hACD2, 16'hB4D3, 16'hBD14, 16'hC556, 16'hB514, 16'h6ACA, 16'h7B4D, 16'hB514, 16'hACD4, 16'hAD15, 16'hBD56, 16'hC597, 16'hC597, 16'hA4D4, 16'h49C6, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hEF1D, 16'hEF5D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8C51, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h7BCF, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8C51, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9CD3, 16'h9492, 16'h9492, 16'h8C51, 16'h9492, 16'h8C51, 16'h9CD3, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'hB596, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFF9E, 16'hF6DB, 16'hEE9A, 16'hF75D, 16'hFF9F, 16'hFFDF, 16'hFF5E, 16'hEE9A, 16'hDDD7, 16'hD555, 16'hCC93, 16'hAB4E, 16'hAB0D, 16'hCC52, 16'hE597, 16'hEDD8, 16'hEE19, 16'hF619, 16'hF65A, 16'hE597, 16'hB38F, 16'hC493, 16'hEE5A, 16'hFEDC, 16'hE659, 16'hDDD7, 16'hDDD7, 16'hE659, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h8BCF, 16'h6289, 16'h51C5, 16'h51C6, 16'h7B0A, 16'h834C, 16'h6207, 16'h6207, 16'h59C6, 16'h838C, 16'h8B8D, 16'h3000, 16'h840F, 16'hC617, 16'hBDD7, 16'hC5D7, 16'hC5D7, 16'hCE18, 16'hD618, 16'h838E, 16'h4943, 16'h93CE, 16'h9C0F, 16'h7B0A, 16'h2800, 16'hB4D2, 16'hD617, 16'hCDD6, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD6, 16'hCDD6, 16'hD5D7, 16'hCDD6, 16'h8BCE, 16'h4080,
        16'hA410, 16'hDE59, 16'hEE9B, 16'hE65A, 16'hDE5A, 16'hDE59, 16'hD659, 16'hCE18, 16'hC5D8, 16'hBD97, 16'hBD96, 16'hC5D7, 16'hCE18, 16'hC618, 16'hC618, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hBDD7, 16'hC5D7, 16'h9451, 16'h6288, 16'h8BCD, 16'h6288, 16'h8BCE, 16'hACD3, 16'h7B4C, 16'h5208, 16'hB4D4, 16'hACD3, 16'h9C51, 16'h8C10, 16'h838F, 16'h8BD0, 16'hAD15, 16'hBD97, 16'h8BCF, 16'h6B0B, 16'hF79D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1D, 16'hCDD9, 16'hC599, 16'hC599, 16'hD65B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8C51, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8C51, 16'h9492, 16'h9CD3, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hF75D, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hEE9A, 16'hC492, 16'hB34F, 16'hAACC, 16'hBBD0, 16'hCC12, 16'hCC53, 16'hD494, 16'hCC52, 16'hB34E, 16'hBB8F, 16'hDD56, 16'hF6DC, 16'hFF9E, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFF9F, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h4100, 16'h7B0B, 16'hB4D3, 16'hB514, 16'hBD14, 16'hC555, 16'hC555, 16'hC555, 16'hBD14, 16'hBD14, 16'hCD96, 16'hA451, 16'h3902, 16'hB595, 16'hC617, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hCE18, 16'hD618, 16'hB514, 16'h4143, 16'h8B8D, 16'h8B8C, 16'h4984, 16'h5A06, 16'hCD95, 16'hCDD7, 16'hCDD6, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD6, 16'hCDD6, 16'hD5D7, 16'hC554, 16'h72CA, 16'h7289, 16'hBD14, 16'hE69A, 16'hE69B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE5A, 16'hD619, 16'hCE18, 16'hCE18, 16'hCE18, 16'hC5D8, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC618, 16'hAD14, 16'h8BCD, 16'hBD14, 16'h8BCF, 16'h7B8D, 16'h6289, 16'h4A07, 16'hACD3, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hA493, 16'h9C52, 16'hBD56, 16'hA493, 16'h41C5, 16'hD659, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD61A, 16'hC5D9, 16'hCDDA, 16'hCDDA, 16'hC599, 16'hE6DD, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hEF5D, 16'h9492, 16'h9492, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8C51, 16'h8C51, 16'hCE59, 16'hDEDB, 16'h8410, 16'h9492, 16'h9492, 16'h8410, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hBDD7, 16'h9492, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hE69A, 16'hDE18, 16'hD596, 16'hDDD8, 16'hE659, 16'hE659, 16'hEE5A, 16'hD515, 16'hB38F, 16'hBB8F, 16'hCC93, 16'hD555, 16'hD556, 16'hDD96, 16'hDDD7, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE99, 16'h59C5, 16'hAC92, 16'hBD54, 16'hBD14, 16'hC555, 16'hC555, 16'hBD55, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD55, 16'hB514, 16'h4145, 16'h83CF, 16'hC617, 16'hBDD7, 16'hC5D7, 16'hC5D7, 16'hCDD8, 16'hCE18, 16'hD618, 16'hCDD7, 16'h6ACA, 16'h6247, 16'h8B4B, 16'h4102, 16'h830B, 16'hCD96, 16'hCDD7, 16'hCDD6, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7,
        16'hCDD7, 16'hCDD6, 16'hCDD6, 16'hCDD7, 16'hCDD6, 16'hCDD7, 16'hD5D7, 16'hAC51, 16'h50C0, 16'h93CE, 16'hE69A, 16'hF71C, 16'hE69B, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hD659, 16'hCE18, 16'hCE18, 16'hC5D8, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC617, 16'hBD96, 16'hC5D7, 16'h9450, 16'hA451, 16'hCDD7, 16'hB514, 16'h62CA, 16'h3984, 16'hACD3, 16'hC596, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD57, 16'hBD57, 16'hBD56, 16'hBD97, 16'h730D, 16'h8C0F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE1A, 16'hC5D9, 16'hCDD9, 16'hCDD9, 16'hC598, 16'hEF1D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9CD3, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h8C51, 16'h8C51, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h9451, 16'h8C51, 16'hDEDB, 16'hFFDF, 16'hEF5D, 16'h9492, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8C51, 16'h8C51, 16'hB596, 16'hFFDF, 16'hE71C, 16'h9492, 16'h8C51, 16'h9CD3, 16'h8410, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h7BCF, 16'h9492, 16'h8410, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hE65A, 16'hDDD7, 16'hDDD7, 16'hDE18, 16'hEEDB, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'h6A48, 16'h6247, 16'h834D, 16'h834D, 16'h93CF, 16'hBCD3, 16'hBD14, 16'hB492, 16'hB4D3, 16'hBD14, 16'hB4D3, 16'hB4D3, 16'h72CB, 16'h3080, 16'hB595, 16'hC617, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hCE18, 16'hCE18, 16'hD618, 16'hD659, 16'hACD3, 16'h38C1, 16'h6A88, 16'h4943, 16'hAC91, 16'hCDD6, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD6, 16'hCDD6, 16'hCDD7, 16'hD617, 16'hCD95, 16'h938D, 16'h2000, 16'hB4D3, 16'hF75D, 16'hFF5D, 16'hF71C, 16'hEEDB, 16'hE69B, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE65A, 16'hE65A, 16'hE69A, 16'hDE59, 16'hCE18, 16'hCE18, 16'hC618, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hA492, 16'hC5D7, 16'h9450, 16'hB4D3, 16'hB514, 16'h5207, 16'h5248, 16'hB515, 16'hC597, 16'hBD56, 16'hBD56,
        16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD57, 16'hACD4, 16'h5208, 16'hAD14, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69C, 16'hC599, 16'hC5D9, 16'hC5D9, 16'hDE9B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8C51, 16'h8C51, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8C51, 16'h8410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8C51, 16'h8C51, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h9492, 16'h8410, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'hA514, 16'hE71C, 16'hFFDF, 16'hDEDB, 16'h8C51,
        16'h9492, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hA514, 16'h8410, 16'h9CD3, 16'h7BCF, 16'hD69A, 16'hFFDF, 16'hD69A, 16'h7BCF, 16'h9492, 16'h8410, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD618, 16'h5943, 16'h8B4D, 16'hAC51, 16'hAC92, 16'hBCD3, 16'hBCD3, 16'hBCD4, 16'hBCD4, 16'hBCD3, 16'h9C10, 16'hA451, 16'hAC92, 16'h6289, 16'h4985, 16'h940F, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hCE18, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'h838D,
        16'h1000, 16'h6248, 16'hCDD6, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD6, 16'hCDD6, 16'hD5D7, 16'hD5D6, 16'hAC92, 16'h5103, 16'h7A89, 16'hDE58, 16'hFFDF, 16'hFF9E, 16'hF71D, 16'hF71C, 16'hEEDC, 16'hEEDB, 16'hE69B, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hD619, 16'hCE18, 16'hCE18, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC618, 16'hAD14, 16'hA491, 16'hC596, 16'h9C50, 16'h9C50, 16'h49C5, 16'h6249, 16'hACD2, 16'hB4D4, 16'hB514, 16'hBD56, 16'hC597, 16'hBD56, 16'hB556, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD57, 16'hA493, 16'h4986, 16'h838E, 16'h8C10, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF75E, 16'hEF5E, 16'hEF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8C51, 16'h8C51, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8C51, 16'h8C51, 16'hB5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h9492, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8C51, 16'h9492, 16'h9492, 16'hDEDB, 16'hEF5D, 16'hAD55, 16'h8410, 16'h8410, 16'hB596, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8C51, 16'h9CD3, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hC618, 16'hA514, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD618, 16'h5080, 16'hA410, 16'hCD55, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hBD14, 16'hBD14, 16'hC555, 16'hAC52, 16'h7B0C, 16'h49C7, 16'h5249, 16'h9C50, 16'hA492, 16'hC617, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hCE17, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hDE59, 16'hC595, 16'h4040, 16'hB4D2, 16'hDE18, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD6, 16'hCDD7, 16'hD617, 16'hCD55, 16'h7B0B, 16'h3000, 16'hAC50, 16'hEF1B, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFF5E, 16'hF71D, 16'hF71C, 16'hEEDC, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69A, 16'hE65A, 16'hE69A, 16'hDE59, 16'hCE18, 16'hCDD8, 16'hCDD7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7,
        16'h940F, 16'hC595, 16'hACD2, 16'h7B0B, 16'h4143, 16'h7B0C, 16'hB492, 16'hA451, 16'h9C10, 16'h93CF, 16'h838E, 16'hA452, 16'hB515, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD97, 16'hACD4, 16'h8BD0, 16'h6ACC, 16'h2802, 16'hB555, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8C51, 16'h8C51, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8C51, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8C51, 16'h9492, 16'h8C51, 16'hD69A, 16'hFFDF, 16'hEF5D,
        16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'h8C51, 16'h8C51, 16'h9CD3, 16'h8410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h7BCF, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE58, 16'h5100, 16'h9C10, 16'hCD55, 16'hC515, 16'hC514, 16'hC514, 16'hC514, 16'hC514, 16'hC514, 16'hC514, 16'hBCD4, 16'hBD14, 16'h49C6, 16'h5248, 16'hBD95, 16'hA491,
        16'hA4D2, 16'hC617, 16'hBDD7, 16'hC5D7, 16'hC5D7, 16'hCE18, 16'hD618, 16'hD619, 16'hD619, 16'hD619, 16'hD659, 16'hE659, 16'hA40F, 16'h834C, 16'hDE18, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hCDD6, 16'hCDD6, 16'hD617, 16'hD5D7, 16'hAC91, 16'h6185, 16'h6985, 16'hD617, 16'hFFDE, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFF5E, 16'hF71D, 16'hF71C, 16'hEEDB, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE65A, 16'hD618, 16'hCE18, 16'hCDD7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC618, 16'hAC92, 16'hB4D2, 16'hBD13, 16'h6207, 16'h4102, 16'h93CF, 16'hC556, 16'hB493, 16'hA3D0, 16'hAC92, 16'hB4D4, 16'hB4D4, 16'h9C52, 16'h9410, 16'h9C51, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD57, 16'hB516, 16'hB556, 16'h9411, 16'h4A08, 16'hB595, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8C51, 16'h8C51, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hAD55, 16'hE71C, 16'hBDD7, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hD69A, 16'h8410, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'h8410, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hCE59, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hCE17, 16'hBD13, 16'h5985, 16'h8B8E, 16'hCD55, 16'hC515, 16'hC515, 16'hC514, 16'hC514, 16'hC514, 16'hC515, 16'hC514, 16'hC514, 16'hC514, 16'hC515, 16'h7B0C, 16'h7B4D, 16'hCDD7, 16'hA491, 16'hAD13, 16'hC618, 16'hBDD7, 16'hC5D7, 16'hC5D7, 16'hCE18, 16'hD618, 16'hD618, 16'hD619, 16'hD659, 16'hDE59, 16'hEE9B, 16'hE659, 16'h7A89, 16'hAC92, 16'hDE18, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hCDD6, 16'hCDD7, 16'hD5D7, 16'hCD55, 16'h8B4D, 16'h2800, 16'h9C10, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFF5E, 16'hFF5D, 16'hF71C, 16'hEEDC, 16'hEEDC, 16'hEEDB, 16'hEEDB, 16'hEE9B,
        16'hE69A, 16'hE65A, 16'hDE59, 16'hD618, 16'hCDD8, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hCE18, 16'hB514, 16'h9BCE, 16'hBCD2, 16'h6A48, 16'h4985, 16'hAC52, 16'hCD56, 16'hC516, 16'hC556, 16'hBD15, 16'hB4D4, 16'h9C10, 16'h93D0, 16'hACD4, 16'hBD56, 16'hA452, 16'h838F, 16'hACD4, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hB556, 16'hB515, 16'hB556, 16'h734D, 16'h5A48, 16'hCE17, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59,
        16'h8410, 16'h9CD3, 16'h8C51, 16'h8410, 16'h8C51, 16'h9492, 16'h8C51, 16'h8C51, 16'h9492, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hB596, 16'h9CD3, 16'h9CD3, 16'hAD55, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h7ACA, 16'h8289, 16'h6185, 16'h9BCF, 16'hCD15, 16'hC515, 16'hC515, 16'hC515,
        16'hC515, 16'hC515, 16'hC515, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hBCD3, 16'hCD55, 16'h9C10, 16'h5207, 16'hC596, 16'hA491, 16'hAD13, 16'hC618, 16'hBDD7, 16'hC5D7, 16'hC618, 16'hCE18, 16'hD618, 16'hD619, 16'hD619, 16'hDE59, 16'hDE59, 16'hE69A, 16'hF6DC, 16'hD596, 16'h5942, 16'hC555, 16'hDE18, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD617, 16'hD5D7, 16'hAC50, 16'h5000, 16'h61C6, 16'hCDD7, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hF75D, 16'hF71C, 16'hF6DC, 16'hEEDB, 16'hE69A, 16'hDE59, 16'hD619, 16'hCE18, 16'hC5D8, 16'hC5D7, 16'hC5D7, 16'hC5D8, 16'hC5D7, 16'hA450, 16'h9BCF, 16'h5185, 16'h72CA, 16'hBD14, 16'hCD97, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hB514, 16'hA451, 16'h8B8E, 16'hB514, 16'hB515, 16'h7B4E, 16'hA453, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD97, 16'hB515, 16'hAD15, 16'h9C93, 16'h628A, 16'h9410, 16'h7B8D, 16'h9451, 16'hDE9A,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9CD3, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hF79E, 16'hE71C, 16'hD69A, 16'hBDD7, 16'hAD55, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8410, 16'h8C51, 16'h9492, 16'h8C51, 16'h8410, 16'hB596, 16'hDEDB, 16'h9CD3, 16'h9CD3, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF75D, 16'hE69A, 16'h61C6, 16'h9BCF, 16'hBC92, 16'hB452, 16'hCD56, 16'hC515, 16'hC515, 16'hCD15, 16'hC515, 16'hB493, 16'hA410, 16'hA410, 16'hAC10, 16'h938E, 16'h9BCF, 16'hA3D0, 16'hC515, 16'hBCD3, 16'h3880, 16'hACD2, 16'hACD2, 16'hAD13, 16'hC618, 16'hC5D7, 16'hC5D7, 16'hCE18, 16'hCE18, 16'hD619, 16'hDE19, 16'hDE59, 16'hDE59, 16'hE65A, 16'hE69A, 16'hF6DC, 16'hFF1D, 16'hAC91, 16'h6A48, 16'hD5D7, 16'hDE18, 16'hDE18, 16'hDE18, 16'hD555, 16'h8ACB, 16'h5080, 16'hBCD3, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hF71D, 16'hF6DC, 16'hE69B, 16'hDE5A, 16'hD619, 16'hCE18, 16'hCDD8, 16'hC5D7, 16'hC5D7, 16'hCDD8, 16'hA450, 16'h938D, 16'h6206, 16'h938E, 16'hCD96, 16'hCD57, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hB4D4, 16'h8B8F, 16'hA492, 16'hBD56, 16'h8B8F, 16'hA493, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD56, 16'hC597, 16'h8C11, 16'h9C93, 16'h9411, 16'h838F, 16'hBD97, 16'hACD4, 16'h734E, 16'h3904, 16'h8C10, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55,
        16'h8C51, 16'h9492, 16'hAD55, 16'hAD55, 16'h9492, 16'h8C51, 16'h8410, 16'h8C51, 16'h8C51, 16'h8C51, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'hAD55, 16'hA514, 16'hAD55, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB,
        16'hAC0F, 16'hA38E, 16'hA3CE, 16'h934E, 16'hC514, 16'hC4D3, 16'hCD15, 16'hC515, 16'hC515, 16'hCD15, 16'hBCD3, 16'h9BCF, 16'h9BCF, 16'hAC10, 16'hAC10, 16'hA410, 16'hBCD3, 16'hC4D4, 16'hC514, 16'hC515, 16'hCD56, 16'h830C, 16'h7B0C, 16'hB4D3, 16'hAD14, 16'hC618, 16'hC5D7, 16'hC5D8, 16'hCE18, 16'hD618, 16'hD619, 16'hDE59, 16'hDE59, 16'hDE59, 16'hE65A, 16'hE65A, 16'hF6DC, 16'hFF5D, 16'hFF1C, 16'h830B, 16'h8B8D, 16'hE659, 16'hDE18, 16'hAC92, 16'h4800, 16'h934C, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hF75D, 16'hEEDB, 16'hE65A, 16'hDE59, 16'hD618, 16'hCE18, 16'hC5D8, 16'hD619, 16'hA492, 16'h7288, 16'h728A, 16'hB492, 16'hD597, 16'hD597, 16'hCD57, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hBD56, 16'hBD56, 16'hC556, 16'hC556, 16'hA451, 16'h9411, 16'hBD55, 16'h9C51, 16'hACD3, 16'hBD56,
        16'hBD56, 16'hBD56, 16'hBD97, 16'hAD15, 16'h734D, 16'hB515, 16'h7B4E, 16'hACD5, 16'hC597, 16'hBD57, 16'hBD57, 16'h9C94, 16'h4A09, 16'h3104, 16'hAD55, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8C51, 16'h9492, 16'h8C51, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'h8C51, 16'h8410, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC555, 16'h828A, 16'hCD15, 16'hE5D7, 16'hAC11, 16'h7209, 16'hBC93, 16'hCD55, 16'hC515, 16'hC514, 16'hC514, 16'hAC11, 16'h9B8F, 16'hBC92, 16'hAC10, 16'h9B8E, 16'hA3D0, 16'hAC51, 16'hBCD4, 16'hC515, 16'hC515, 16'hC515, 16'hCD55, 16'hB493, 16'h4985, 16'h938E, 16'hACD3, 16'hCE18, 16'hC5D7, 16'hCDD8, 16'hCE18, 16'hD618, 16'hD619, 16'hDE59, 16'hDE59, 16'hE65A, 16'hE65A, 16'hE69A, 16'hF6DC, 16'hFF1D, 16'hFF9E, 16'hEE9A, 16'h7207, 16'hA450, 16'h93CE, 16'h5903,
        16'hC555, 16'hFF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hE69B, 16'hE65A, 16'hD619, 16'hD619, 16'hD618, 16'hAC51, 16'h5902, 16'h82CB, 16'hAC11, 16'hB452, 16'hAC11, 16'hB493, 16'hCD56, 16'hCD57, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hBD56, 16'hC556, 16'hBD16, 16'hBD16, 16'hC556, 16'hA453, 16'h93D0, 16'hB515, 16'h93D0, 16'hB515, 16'hBD97, 16'hBD56, 16'hBD97, 16'h83D0, 16'h9C92, 16'h9451, 16'h9C52, 16'hC598, 16'hBD57, 16'hBD57, 16'hBD57, 16'hBD98, 16'hB557, 16'h9453, 16'h62CB, 16'h7B8E, 16'hAD55, 16'hF79D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h7BCF, 16'h8C51, 16'h8410, 16'h8C51, 16'h9492, 16'h9CD3, 16'hAD55, 16'hC618, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hA410, 16'h9B8F, 16'hE619, 16'hF69B, 16'hDD98, 16'hCD15, 16'h7A49, 16'h9B8F, 16'hCD55, 16'hC515, 16'hC514, 16'hA3D0, 16'hA3CF, 16'hB452, 16'h9B4E, 16'h9B8E, 16'hBC93, 16'hC515, 16'hCD15, 16'hCD15, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hCD55, 16'h830C, 16'h6A08, 16'hB4D3, 16'hCE18, 16'hCDD7, 16'hCE18, 16'hCE18, 16'hD618, 16'hDE59, 16'hDE59, 16'hDE59, 16'hE69A, 16'hE69A, 16'hE69A, 16'hF6DC, 16'hFF5D, 16'hFF5E, 16'hFEDC, 16'h9B8D, 16'h3000, 16'h5000, 16'hC514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hF71C, 16'hE69B, 16'hE69A, 16'hD618, 16'h8B8D, 16'h5000, 16'hC4D3, 16'hE597, 16'hC4D4, 16'hB452, 16'hA3D0, 16'hAC11, 16'h9B8E, 16'hC4D4, 16'hD597, 16'hC556, 16'hCD56, 16'hC556,
        16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hBD16, 16'hBD16, 16'hC557, 16'h9C52, 16'h9411, 16'hB514, 16'h8C10, 16'hBD56, 16'hBD97, 16'hA492, 16'h9C52, 16'hA493, 16'h83CF, 16'hC597, 16'hC557, 16'hBD57, 16'hBD97, 16'hBD97, 16'hBD57, 16'hBD57, 16'hBD98, 16'hB557, 16'h9452, 16'h3986, 16'h734C, 16'hCE58, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'hB596, 16'hCE59, 16'hDEDB, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'h934C, 16'hC4D4, 16'hF6DC, 16'hFE9C, 16'hEE19, 16'hE5D9, 16'hE5D8, 16'hB452, 16'h9B4D, 16'hCD15, 16'hCD15, 16'hA3CF, 16'hA410, 16'hAC11, 16'h8B0D, 16'hBC92, 16'hCD15, 16'hCD15, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hCD55, 16'hD556, 16'hC514, 16'h5986, 16'h9BCF, 16'hD618, 16'hCDD8, 16'hCE18, 16'hD618, 16'hD619, 16'hDE59, 16'hDE59,
        16'hE69A, 16'hE69A, 16'hE69B, 16'hEE9B, 16'hF6DC, 16'hFF5E, 16'hD5D7, 16'h7A09, 16'h7248, 16'h6A07, 16'h9BCE, 16'h930C, 16'hD596, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hF71D, 16'hD5D7, 16'h6A07, 16'h7208, 16'hDD96, 16'hF65A, 16'hF61A, 16'hEDD9, 16'hD557, 16'hBC93, 16'hB452, 16'hC4D4, 16'hA3D0, 16'hBC93, 16'hD597, 16'hCD56, 16'hCD57, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hBD56, 16'hC556, 16'h8BCF, 16'hA493, 16'h9411, 16'hACD4, 16'hB515, 16'h93D0, 16'hACD3, 16'h9452, 16'hBD56, 16'hC597, 16'hBD57, 16'hC557, 16'hC597, 16'hC597, 16'hBD97, 16'hBD57, 16'hBD97, 16'hBD98, 16'hBD98, 16'hAD15, 16'h734E, 16'h2000, 16'h9451, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE18, 16'h9B4C, 16'hE659, 16'hFF5F, 16'hFEDD, 16'hF65A, 16'hEE19, 16'hE5D8, 16'hDD98, 16'hD556, 16'h930D, 16'hBC92, 16'hB452, 16'hA3D0, 16'hB452, 16'h930D, 16'hC4D4, 16'hCD15, 16'hC514, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hCD15, 16'hCD55, 16'hCD15, 16'hBC93, 16'hB492, 16'hDD97, 16'hB452, 16'h2800, 16'hB4D3, 16'hD618, 16'hD618, 16'hD619, 16'hDE59, 16'hDE59, 16'hE65A, 16'hE69A, 16'hEE9B, 16'hEE9B, 16'hEEDB, 16'hFF1D, 16'hEE5A, 16'h8B4C, 16'h8B8E, 16'hA451, 16'hA450, 16'hCD55, 16'hBD13, 16'h6840, 16'hD618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5D, 16'hB493, 16'h7185, 16'hB411, 16'hF619, 16'hF65B,
        16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE5D9, 16'hDDD8, 16'hD556, 16'hB452, 16'hBC93, 16'hA411, 16'hB493, 16'hD597, 16'hCD57, 16'hCD57, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hBD56, 16'hC556, 16'hACD4, 16'h8BD0, 16'hACD4, 16'h9C52, 16'hBD56, 16'hB515, 16'h9411, 16'hB515, 16'hC597, 16'hBD57, 16'hC557, 16'hC557, 16'hC557, 16'hC597, 16'hBD97, 16'hBD97, 16'hBD97, 16'hBD97, 16'hBD97, 16'hBD98, 16'hBD97, 16'h9C53, 16'h41C8, 16'h83CE, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDDD7, 16'h9B4D, 16'hE69A, 16'hFF9F, 16'hFF1D, 16'hF69C, 16'hF65A, 16'hEE19, 16'hE5D8, 16'hDD98, 16'hDD97, 16'hB452, 16'h934D, 16'hBC93, 16'hB452, 16'h9B4E, 16'hC4D4, 16'hCD15, 16'hC514, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hCD15, 16'hC514, 16'hB451, 16'hABD0,
        16'hB451, 16'hB492, 16'hD596, 16'hDD97, 16'h9B8F, 16'h2000, 16'hBD14, 16'hE65A, 16'hDE59, 16'hDE59, 16'hE65A, 16'hE69A, 16'hEEDB, 16'hEEDB, 16'hEEDB, 16'hEEDC, 16'hFF1D, 16'hA410, 16'h93CE, 16'hD617, 16'hD617, 16'hC554, 16'h8B8D, 16'hAC91, 16'hA450, 16'h8ACB, 16'hFF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hA3D0, 16'h8209, 16'hDD56, 16'hFE5B, 16'hF65B, 16'hF65A, 16'hF61A, 16'hF61A, 16'hF65A, 16'hEE1A, 16'hE5D8, 16'hDDD8, 16'hD597, 16'hB452, 16'hBCD4, 16'hAC10, 16'hB493, 16'hCD97, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD57, 16'hC557, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hBD15, 16'h9C11, 16'hB515, 16'hB515, 16'hBD56, 16'hA453, 16'hB515, 16'hC597, 16'hC557, 16'hC557, 16'hC557, 16'hC557, 16'hC557, 16'hC597, 16'hBD97, 16'hBD97, 16'hBD97, 16'hBD97, 16'hBD97, 16'hBD97, 16'hBD97, 16'hBD98, 16'hB516,
        16'h730E, 16'h4A08, 16'hB595, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD55, 16'hB410, 16'hF6DC, 16'hFFDF, 16'hFF5E, 16'hFEDD, 16'hF69B, 16'hEE5A, 16'hE619, 16'hE5D8, 16'hDD98, 16'hDD97, 16'hD556, 16'h9B4E, 16'hBC92, 16'hB451, 16'hC4D3, 16'hCD15, 16'hC514, 16'hC515, 16'hCD15, 16'hCD15, 16'hC515, 16'hCD15, 16'hB493, 16'h9B4E, 16'hB410, 16'hBC93, 16'hAC51, 16'hA3D0, 16'hB451, 16'hDDD8, 16'hDDD7, 16'h82CB, 16'h5945, 16'hDDD7, 16'hE69A, 16'hE65A, 16'hE69A, 16'hEEDB, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hFF1D, 16'hD5D7, 16'h830B, 16'hCE16, 16'hCE17, 16'hCDD6, 16'hCE17, 16'hD5D6, 16'h9C50, 16'h93CE, 16'h7A8A, 16'hCD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hBCD3, 16'h7186, 16'hABD0, 16'hEE19, 16'hFE5B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hF61A, 16'hF65A, 16'hF65A, 16'hEE19, 16'hDD98, 16'hDD98, 16'hDD98, 16'hB452, 16'hBC93, 16'hA3D0, 16'hC515, 16'hCD97, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD57, 16'hC556, 16'hC556, 16'hC556, 16'hBD56, 16'hC556, 16'hA492, 16'hB4D4, 16'hBD56, 16'hBD15, 16'hBD56, 16'hC597, 16'hC597, 16'hC597, 16'hC557, 16'hC557, 16'hC557, 16'hC557, 16'hC557, 16'hBD97, 16'hBD97, 16'hBD97, 16'hBD97, 16'hBD97, 16'hBD97, 16'hBD97, 16'hBD57, 16'hBD98, 16'hBD97, 16'h9C93, 16'h62CB, 16'h9451, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hC4D3, 16'hBC51, 16'hFF5D, 16'hFFDF, 16'hFF9E, 16'hFF1D, 16'hFEDC, 16'hF69B, 16'hEE1A, 16'hE5D9, 16'hDDD8, 16'hDD98, 16'hDD97, 16'hDD97, 16'hBC52, 16'hABD0, 16'hB452,
        16'hCCD4, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC515, 16'hCD55, 16'hAC11, 16'h9B4D, 16'hBC51, 16'hA3CF, 16'h934E, 16'hB452, 16'hCD15, 16'hDD97, 16'hDD97, 16'hDDD8, 16'hDD97, 16'h930D, 16'h6A07, 16'hDDD7, 16'hF6DB, 16'hEE9B, 16'hF6DC, 16'hF71C, 16'hF71C, 16'hF71C, 16'hFF1D, 16'h8B4D, 16'hACD2, 16'hD617, 16'hCDD6, 16'hD617, 16'hD617, 16'hD617, 16'hD657, 16'h9C0F, 16'h7ACA, 16'h7207, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD617, 16'h8A8A, 16'h928B, 16'hE598, 16'hEE1A, 16'hDD56, 16'hEE1A, 16'hF65B, 16'hF65A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hE5D9, 16'hDD98, 16'hDD98, 16'hD597, 16'hAC11, 16'hBC93, 16'h9B8F, 16'hC516, 16'hCD97, 16'hCD57, 16'hCD57, 16'hCD57, 16'hC556, 16'hC556, 16'hBD56, 16'hCD97, 16'hAC93, 16'h8B8F, 16'hBD15, 16'hBD56, 16'hC556, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597,
        16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hBD97, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD98, 16'hB516, 16'h7B8E, 16'h62CA, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hBC92, 16'hC4D4, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hFEDD, 16'hFE9C, 16'hF65A, 16'hEE19, 16'hE5D9, 16'hE5D8, 16'hDDD8, 16'hDD97, 16'hDD97, 16'hCD15, 16'hABD0, 16'hC4D4, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC515, 16'hCD55, 16'hB451, 16'h9B8E, 16'hB451, 16'h9B4D, 16'hB452, 16'hDD56, 16'hE5D8, 16'hE598, 16'hDD98, 16'hDD98, 16'hE5D9, 16'hEE1A, 16'hEDD9, 16'h930C, 16'h6186, 16'hCD96, 16'hF6DC, 16'hF6DC, 16'hF71C, 16'hF71D, 16'hFF5E, 16'hD596, 16'h7B0B, 16'hD617, 16'hCE16, 16'hCE17, 16'hBD54, 16'h940F, 16'hA491, 16'hCDD6, 16'hCDD6, 16'h93CE, 16'h7A89, 16'hBCD2, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'h8B0C, 16'h6800, 16'hBC92, 16'hF619, 16'hCC93, 16'hE598, 16'hED98, 16'hCC94, 16'hEE19, 16'hF65B, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF65A, 16'hEE1A, 16'hDD98, 16'hDD98, 16'hDD98, 16'hCD15, 16'hAC11, 16'hB452, 16'hAC11, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD57, 16'hC556, 16'hC556, 16'hCD56, 16'hA451, 16'h9B8F, 16'hC515, 16'hC557, 16'hC557, 16'hCD97, 16'hCD97, 16'hCD97, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hBD97, 16'hBD97, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD98, 16'hC598, 16'hBD97, 16'h8BD0, 16'h5208, 16'hC5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hC4D3, 16'hC514, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF5E,
        16'hFEDD, 16'hF69B, 16'hF65A, 16'hEE1A, 16'hEE19, 16'hE5D9, 16'hDD97, 16'hDD97, 16'hDD97, 16'hDD97, 16'hBC52, 16'hB452, 16'hCD15, 16'hCD15, 16'hCD15, 16'hC515, 16'hCD55, 16'hAC10, 16'h9B8E, 16'hAC10, 16'h934D, 16'hCD15, 16'hDD97, 16'hD557, 16'hDD97, 16'hDD97, 16'hE5D8, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hED98, 16'h9B4E, 16'h4000, 16'hBCD3, 16'hF6DB, 16'hFF5E, 16'hFF5E, 16'hFF5D, 16'h830B, 16'hAC91, 16'hD617, 16'hCDD6, 16'hCDD6, 16'h838D, 16'hACD3, 16'hA450, 16'h834C, 16'hD617, 16'h9C0F, 16'h9BCF, 16'h7A08, 16'hD5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD618, 16'h934D, 16'h7144, 16'hB411, 16'hEDD9, 16'hFE5B, 16'hF65B, 16'hDD57, 16'hBBD1, 16'hE557, 16'hF619, 16'hD4D5, 16'hF61A, 16'hF65B, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hE5D9, 16'hDD98, 16'hDD98, 16'hDD98, 16'hB453, 16'hB452, 16'hAC11, 16'hBCD4, 16'hD597, 16'hCD57, 16'hCD56, 16'hCD57, 16'hD556, 16'h9BCF,
        16'h938F, 16'hCD56, 16'hD597, 16'hCD97, 16'hD5D8, 16'hD5D8, 16'hCD97, 16'hCD97, 16'hCD97, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hBD97, 16'hBD97, 16'hBD97, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD97, 16'hBD98, 16'hBD98, 16'h9C53, 16'h3905, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hC514, 16'hCD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF1E, 16'hF69C, 16'hF65B, 16'hEE5A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hDDD8, 16'hDD97, 16'hDD97, 16'hDD97, 16'hD556, 16'hAC11, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD56, 16'hBC93, 16'hA38E, 16'hABCF, 16'h9B8E, 16'hCD55, 16'hD557, 16'hD556, 16'hD557, 16'hDD97, 16'hEDD9, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hF61A, 16'hE557, 16'hE5D8, 16'hEE1A, 16'hB452, 16'h5000, 16'h8ACB, 16'hE618, 16'hFF5E, 16'hEE9A, 16'h5903, 16'hC554, 16'hD616, 16'hD617, 16'hBD54,
        16'hA491, 16'hD617, 16'hDE17, 16'h9C10, 16'hACD2, 16'hAC91, 16'hAC51, 16'hAC51, 16'h6103, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hCD96, 16'h934C, 16'h79C7, 16'hC493, 16'hEDD9, 16'hFE5B, 16'hF65B, 16'hF65A, 16'hF61A, 16'hF65B, 16'hF61A, 16'hC453, 16'hE598, 16'hED98, 16'hCCD4, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hEE1A, 16'hE5D9, 16'hDD98, 16'hDD98, 16'hD557, 16'hA3D0, 16'hB452, 16'h9B8F, 16'hCD56, 16'hCD56, 16'hD597, 16'hCD55, 16'h934E, 16'hAC10, 16'hD596, 16'hD597, 16'hD597, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hD597, 16'hCD97, 16'hCD97, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hBD97, 16'hBD97, 16'hBD97, 16'hBD97, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD98, 16'hA493, 16'h4104, 16'hBDD6, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC514, 16'hCD14, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hFEDC, 16'hF69B, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hE5D9, 16'hDDD8, 16'hDD98, 16'hDD97, 16'hDD97, 16'hCD15, 16'hBC93, 16'hD556, 16'hCD15, 16'hCD15, 16'hA38F, 16'hB410, 16'hABCF, 16'hD556, 16'hD556, 16'hCD56, 16'hD556, 16'hDD97, 16'hEE19, 16'hEE1A, 16'hEE19, 16'hF61A, 16'hEE19, 16'hCCD4, 16'hCC94, 16'hF61A, 16'hEE1A, 16'hF61A, 16'hDD57, 16'h9B0D, 16'h5800, 16'hA3CF, 16'hAC51, 16'h934D, 16'hD5D7, 16'hD617, 16'hD617, 16'hB513, 16'h9C50, 16'hD5D6, 16'hD5D7, 16'hAC92, 16'h9C10, 16'hB4D3, 16'hA410, 16'hE618, 16'h6A08, 16'hC596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hCDD7, 16'h9C10, 16'h8A89, 16'hA34D, 16'hCCD4, 16'hEE19, 16'hFE5B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65B, 16'hF65B, 16'hF61A, 16'hF65B, 16'hEDD9, 16'hC411, 16'hF5D9, 16'hD4D5, 16'hDD56, 16'hF65B, 16'hEE1A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hEE1A,
        16'hDD98, 16'hDD98, 16'hDD98, 16'hBC93, 16'hABD0, 16'hA38F, 16'hC4D4, 16'hD597, 16'hC514, 16'h934E, 16'hB492, 16'hDD97, 16'hD597, 16'hD597, 16'hE5D9, 16'hEE1A, 16'hE619, 16'hE619, 16'hDDD9, 16'hD5D8, 16'hCD97, 16'hCD97, 16'hCD97, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hBD97, 16'hBD97, 16'hBD97, 16'hBD97, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD98, 16'hA494, 16'h4986, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD55, 16'hCD14, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hFEDD, 16'hFEDC, 16'hF65B, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hE5D9, 16'hE5D8, 16'hDDD8, 16'hDD98, 16'hDD97, 16'hD557, 16'hC493, 16'hC515, 16'hD556, 16'hBC92, 16'hA38E, 16'hA38E, 16'hCD15, 16'hD556, 16'hCD56, 16'hD556, 16'hD597, 16'hEDD9, 16'hEE19, 16'hEE19, 16'hF61A, 16'hDD56, 16'hD515, 16'hBC11, 16'hF61A, 16'hEE1A,
        16'hEE1A, 16'hEE1A, 16'hF65B, 16'hF65A, 16'hD515, 16'h8ACC, 16'h4000, 16'h69C7, 16'hA40F, 16'hBD13, 16'hD5D6, 16'hCD96, 16'hA450, 16'hD5D7, 16'hDE18, 16'hA491, 16'hA492, 16'hBD14, 16'h9BCF, 16'hEE9A, 16'hBD13, 16'h9B8E, 16'hFF5E, 16'hFFDF, 16'hF75D, 16'hDE9A, 16'hB514, 16'h834C, 16'h7207, 16'h8249, 16'hB451, 16'hE597, 16'hF65A, 16'hF69B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hFE5B, 16'hDD16, 16'hCC93, 16'hF5D9, 16'hCC93, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hE5D9, 16'hDD97, 16'hDD98, 16'hD557, 16'hB411, 16'hAC11, 16'hCD14, 16'hC4D4, 16'h930D, 16'hC4D4, 16'hDDD8, 16'hD597, 16'hD597, 16'hE5D9, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hDDD8, 16'hD598, 16'hCD97, 16'hCD97, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hBD97, 16'hBD97, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD97, 16'hC5D8,
        16'hA493, 16'h51C7, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD597, 16'hCD14, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hFF1D, 16'hFEDC, 16'hFEDC, 16'hFE9C, 16'hF65B, 16'hF65A, 16'hF65A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hE5D8, 16'hDD98, 16'hDD98, 16'hD556, 16'hB452, 16'hD515, 16'hABCF, 16'hBC10, 16'hBC93, 16'hD597, 16'hD556, 16'hD556, 16'hD557, 16'hE5D9, 16'hEE1A, 16'hEE19, 16'hF61A, 16'hDD15, 16'hD4D4, 16'hC452, 16'hEE1A, 16'hEE1A, 16'hF61A, 16'hF65A, 16'hF65A, 16'hEE1A, 16'hEE5A, 16'hF65B, 16'hF65A, 16'hDD56, 16'hABD0, 16'h7208, 16'h5080, 16'h7A89, 16'h9BCF, 16'h9BCE, 16'hAC91, 16'hC554, 16'hA40F, 16'hBD14, 16'hC554, 16'h9BCF, 16'hE5D7, 16'hBCD2, 16'h8ACB, 16'hB451, 16'h934E, 16'h7248, 16'h6040, 16'h8249, 16'hB451, 16'hD555, 16'hEDD8, 16'hFE5B, 16'hF65B, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A,
        16'hF65A, 16'hCC52, 16'hE598, 16'hDD16, 16'hDD16, 16'hF65B, 16'hF61A, 16'hF61A, 16'hF61A, 16'hEE1A, 16'hEE5A, 16'hF65A, 16'hEE19, 16'hDD97, 16'hDD97, 16'hDD97, 16'hD557, 16'hB411, 16'hAC10, 16'hA38F, 16'hCD16, 16'hDDD8, 16'hD597, 16'hDD98, 16'hE619, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE61A, 16'hE5D9, 16'hD5D8, 16'hCD98, 16'hCD97, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hBD97, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD97, 16'hC5D8, 16'h9C52, 16'h6A8B, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE19, 16'hCD14, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hFF1D, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hF65B, 16'hF65B, 16'hF65A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hE598, 16'hE5D8, 16'hC493, 16'hBC51, 16'hC451, 16'hB3CF, 16'hCD15, 16'hD597, 16'hD556,
        16'hD557, 16'hE5D9, 16'hEE1A, 16'hEDD9, 16'hEE1A, 16'hE557, 16'hBC10, 16'hCC93, 16'hDD56, 16'hF65B, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE1A, 16'hEE1A, 16'hF65A, 16'hF65A, 16'hEDD8, 16'hDD56, 16'hBC92, 16'h9B4D, 16'h824A, 16'h71C6, 16'h6142, 16'h50C0, 16'h7A89, 16'h82CA, 16'h5943, 16'h7A07, 16'h71C7, 16'h8ACC, 16'h930C, 16'hBC52, 16'hD556, 16'hE5D8, 16'hF65A, 16'hFE9B, 16'hED98, 16'hC452, 16'hE597, 16'hDD56, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hFE5B, 16'hE557, 16'hCC93, 16'hF5D9, 16'hCC53, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hE5D9, 16'hDD97, 16'hDD97, 16'hDD98, 16'hDD97, 16'hA3CF, 16'hAC10, 16'hDD97, 16'hE5D8, 16'hDD98, 16'hE5D8, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hDDD8, 16'hD598, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD98, 16'hCD97, 16'hCD97, 16'hC597, 16'hC597,
        16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC598, 16'hC598, 16'hC598, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD98, 16'hBD98, 16'hC5D8, 16'h9411, 16'h7B4D, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hC492, 16'hFF1D, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hFEDC, 16'hFE9C, 16'hFEDC, 16'hFEDC, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9B, 16'hF65B, 16'hF65A, 16'hEE1A, 16'hEE19, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D8, 16'hB410, 16'hD4D4, 16'hCCD3, 16'hDD97, 16'hDD97, 16'hDD97, 16'hE5D8, 16'hEE1A, 16'hEE19, 16'hEE1A, 16'hEDD9, 16'hC452, 16'hDD15, 16'hD515, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hF65A, 16'hD515, 16'hDD15, 16'hE597, 16'hFE5B, 16'hF61A, 16'hEE1A, 16'hE598, 16'hDD57, 16'hCD15, 16'hCD15, 16'hC493, 16'hBC93, 16'hD515, 16'hE597, 16'hEE1A, 16'hF61A, 16'hFE5B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hEE1A, 16'hF61B, 16'hDD16, 16'hDD15, 16'hD4D5,
        16'hE5D8, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hF65A, 16'hC453, 16'hED98, 16'hD494, 16'hE598, 16'hF65A, 16'hEE1A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hE5D8, 16'hDD98, 16'hDDD8, 16'hD515, 16'h9B4E, 16'hBC93, 16'hE5D8, 16'hDD98, 16'hE5D8, 16'hEE19, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hDDD9, 16'hDDD8, 16'hD598, 16'hD5D8, 16'hDDD8, 16'hDDD9, 16'hE5D9, 16'hDDD9, 16'hDDD9, 16'hDDD8, 16'hD598, 16'hD598, 16'hCD97, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC598, 16'hBD98, 16'hC598, 16'hBD98, 16'hBD98, 16'hBD98, 16'hC597, 16'h730C, 16'hA4D3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hBC51, 16'hEE5A, 16'hFFDF, 16'hFF9E, 16'hFF1D, 16'hFEDC, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9B, 16'hF65B, 16'hEE1A, 16'hEE19, 16'hEE19,
        16'hE619, 16'hE5D9, 16'hE619, 16'hEE19, 16'hEE19, 16'hEE19, 16'hDD56, 16'hB3D0, 16'hDD97, 16'hDDD8, 16'hDD97, 16'hE5D8, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE1A, 16'hD515, 16'hDD15, 16'hD4D4, 16'hE598, 16'hF65A, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hDD56, 16'hBC11, 16'hDCD5, 16'hDD15, 16'hF61A, 16'hEE1A, 16'hF65A, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hFE5B, 16'hFE5B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61B, 16'hF61A, 16'hD4D4, 16'hDD56, 16'hD516, 16'hF65B, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hF65B, 16'hDD56, 16'hD4D5, 16'hE556, 16'hD516, 16'hF65B, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hE619, 16'hE5D9, 16'hDDD8, 16'hBC93, 16'h9B0D, 16'hCCD5, 16'hE5D9, 16'hE5D9, 16'hEE19, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A,
        16'hE61A, 16'hE619, 16'hE619, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE619, 16'hE5D9, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD8, 16'hD5D8, 16'hD598, 16'hCD98, 16'hCD97, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC598, 16'hC598, 16'hC598, 16'hC598, 16'hBD97, 16'hC5D8, 16'hBD56, 16'h5A07, 16'hCDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBC93, 16'hDDD8, 16'hFF9F, 16'hFF5E, 16'hFF1D, 16'hFEDC, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9B, 16'hFE9B, 16'hF65B, 16'hF65A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hF65A, 16'hD515, 16'hB411, 16'hE5D8, 16'hE5D9, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEDD9, 16'hC452, 16'hE556, 16'hCC93, 16'hF65A, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hC452, 16'hDD16, 16'hD4D4, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hE597, 16'hEDD9, 16'hF61A,
        16'hF61A, 16'hF61A, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hF61A, 16'hFE5B, 16'hD4D4, 16'hDD56, 16'hD4D4, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hCC53, 16'hE557, 16'hCC93, 16'hF61A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hE5D8, 16'hBC52, 16'hBC52, 16'hDD97, 16'hE5D9, 16'hE5D9, 16'hF61A, 16'hF65A, 16'hEE5A, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE5D9, 16'hDDD9, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD9, 16'hD5D8, 16'hD598, 16'hCD98, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC598, 16'hC597, 16'hC598, 16'hC598, 16'hC598, 16'hBD97, 16'hC5D8, 16'hA493, 16'h6A48, 16'hE71B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD55, 16'hCD15, 16'hFF9F, 16'hFF9F, 16'hFF1D, 16'hFEDC, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C,
        16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hF69B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hF61A, 16'hD515, 16'hD515, 16'hEE1A, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hF65A, 16'hD515, 16'hD4D5, 16'hD4D5, 16'hE597, 16'hF65B, 16'hEE1A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hD515, 16'hCC94, 16'hDD16, 16'hE557, 16'hF65B, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hEE19, 16'hC453, 16'hD515, 16'hF61A, 16'hF65A, 16'hF61A, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hF65B, 16'hE556, 16'hD4D5, 16'hDD56, 16'hDD57, 16'hF65B, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF65B, 16'hD4D5, 16'hDD16, 16'hD4D4, 16'hED98, 16'hF65A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hDD57, 16'hD515, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE5A,
        16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hDDD9, 16'hE5D9, 16'hDDD9, 16'hDDD8, 16'hDDD9, 16'hDDD9, 16'hDDD8, 16'hDDD8, 16'hD598, 16'hCD97, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC598, 16'hC598, 16'hC598, 16'hC598, 16'hBD98, 16'hCDD8, 16'h93CF, 16'h834D, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65A, 16'hBC51, 16'hF75D, 16'hFFDF, 16'hFF1D, 16'hFEDC, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hF69B, 16'hFE9B, 16'hF69B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hF61A, 16'hCCD4, 16'hE598, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hCC94, 16'hE557, 16'hCC94, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hD515, 16'hDD15, 16'hD4D4,
        16'hF61A, 16'hEE1A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF65B, 16'hE557, 16'hCC94, 16'hD515, 16'hEE19, 16'hF65A, 16'hF61A, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEDD9, 16'hCC53, 16'hE557, 16'hD4D5, 16'hF65B, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF65B, 16'hE597, 16'hCC93, 16'hDCD5, 16'hDD16, 16'hF65B, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE619, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD8, 16'hDDD8, 16'hD5D8, 16'hCD97, 16'hC597, 16'hC598, 16'hC598, 16'hC598, 16'hC598, 16'hC598, 16'hC598, 16'hC598, 16'hC598, 16'hC556, 16'h6A48, 16'hCE17,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D,
        16'hB3CF, 16'hEE9A, 16'hFFDF, 16'hFF9E, 16'hFF1D, 16'hFEDC, 16'hFEDC, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hEE19, 16'hD4D4, 16'hE598, 16'hF65A, 16'hF61A, 16'hEDD8, 16'hCC94, 16'hDD56, 16'hCCD4, 16'hF65B, 16'hEE1A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hE598, 16'hD515, 16'hE557, 16'hD515, 16'hF65B, 16'hEE1A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF65B, 16'hD515, 16'hD515, 16'hD4D4, 16'hF61A, 16'hF65A, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hF65B, 16'hCC93, 16'hE597, 16'hD4D4, 16'hEE1A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hF5D9, 16'hD4D5, 16'hE557, 16'hD4D4, 16'hF61A,
        16'hEE1A, 16'hF61A, 16'hF61A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hF61A, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hE619, 16'hE5D9, 16'hDDD9, 16'hE5D9, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD8, 16'hD5D8, 16'hD5D8, 16'hCDD8, 16'hC598, 16'hC597, 16'hC598, 16'hC598, 16'hC598, 16'hC598, 16'hC598, 16'hC597, 16'hCDD8, 16'hACD3, 16'h7ACB, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC4D4, 16'hCD55, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hF69B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hEE1A, 16'hF65A, 16'hEDD8, 16'hC493, 16'hE5D9, 16'hF65B, 16'hDD56, 16'hDD16, 16'hD4D5, 16'hDD57, 16'hF65B, 16'hEE1A,
        16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hF65B, 16'hCC94, 16'hE556, 16'hDD16, 16'hEDD8, 16'hF65A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF65A, 16'hCCD4, 16'hDD56, 16'hD4D4, 16'hF61A, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hFE5B, 16'hD4D5, 16'hE557, 16'hD4D4, 16'hDD56, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hEE1A, 16'hF65A, 16'hEDD9, 16'hC452, 16'hEDD9, 16'hF61A, 16'hF61A, 16'hF61A, 16'hEE1A, 16'hEE5A, 16'hEE1A, 16'hF61A, 16'hEE1A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hE61A, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hDDD9, 16'hDDD9, 16'hDDD8, 16'hDDD8, 16'hD5D8,
        16'hD5D8, 16'hD5D8, 16'hCD97, 16'hC598, 16'hC598, 16'hC598, 16'hC598, 16'hC598, 16'hC598, 16'hC598, 16'hC598, 16'h834D, 16'hACD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE18, 16'hBC52, 16'hFF9E, 16'hFFDF, 16'hFF5E, 16'hFEDD, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hEDD8, 16'hCC94, 16'hF619, 16'hE5D8, 16'hEDD9, 16'hD4D4, 16'hE598, 16'hF65B, 16'hEE1A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hC452, 16'hE598, 16'hD4D4, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hEE1A, 16'hF65A, 16'hCCD4, 16'hE557, 16'hCC93, 16'hF61A, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hE557, 16'hDD15, 16'hDD56, 16'hD515, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A,
        16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hEDD9, 16'hCC93, 16'hE557, 16'hF65B, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE5D9, 16'hE5D9, 16'hDDD9, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hD5D8, 16'hDDD8, 16'hD598, 16'hC597, 16'hC597, 16'hC598, 16'hC598, 16'hC598, 16'hC598, 16'hC597, 16'hC598, 16'hB515, 16'h6A89, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hB3CF, 16'hF71C, 16'hFFDF, 16'hFF9F, 16'hFEDD, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A,
        16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hEDD9, 16'hCC93, 16'hDD57, 16'hF65B, 16'hCCD4, 16'hE597, 16'hF65B, 16'hEE1A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE1A, 16'hF65A, 16'hE598, 16'hC452, 16'hE597, 16'hD4D5, 16'hF65B, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hEE1A, 16'hF65A, 16'hCC93, 16'hDD56, 16'hCC93, 16'hF61A, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hEDD8, 16'hD494, 16'hE598, 16'hCCD4, 16'hF65B, 16'hEE1A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hEE1A, 16'hDD56, 16'hC453, 16'hE598, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A,
        16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE5D9, 16'hE5D9, 16'hDDD8, 16'hDDD8, 16'hDDD9, 16'hDDD8, 16'hDDD8, 16'hD5D8, 16'hD598, 16'hC597, 16'hC597, 16'hC598, 16'hC598, 16'hC598, 16'hC598, 16'hC597, 16'hCDD8, 16'h9410, 16'hA450, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC4D3, 16'hD5D7, 16'hFFDF, 16'hFFDF, 16'hFF1E, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9B, 16'hFE9B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hF65B, 16'hEDD9, 16'hEDD8, 16'hE598, 16'hD4D5, 16'hEDD9, 16'hF65A, 16'hEE1A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE1A, 16'hF65B, 16'hDD56, 16'hCC94, 16'hE557, 16'hDD16, 16'hF65B, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hEE1A, 16'hF65A, 16'hCCD4, 16'hE557, 16'hD4D4, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A,
        16'hF65A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hCC93, 16'hE598, 16'hC453, 16'hF61A, 16'hEE1A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hEE19, 16'hDD57, 16'hCC94, 16'hD515, 16'hEDD9, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE619, 16'hE5D9, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hD5D8, 16'hCD98, 16'hC597, 16'hC597, 16'hC598, 16'hC598, 16'hC598, 16'hC597, 16'hC598, 16'hBD56, 16'h7ACB, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE618, 16'hBC51, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFEDC, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hF65B, 16'hEE19, 16'hFE9C, 16'hFE9B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A,
        16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hEDD9, 16'hD515, 16'hE597, 16'hF61A, 16'hF65B, 16'hEE5A, 16'hEE1A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hEE1A, 16'hF65B, 16'hDD56, 16'hD4D5, 16'hDD15, 16'hDD57, 16'hF65B, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hEE1A, 16'hF65A, 16'hCCD4, 16'hE557, 16'hD4D4, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hCC93, 16'hE598, 16'hC493, 16'hEDD9, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE19, 16'hD515, 16'hCC93, 16'hD515, 16'hEDD9, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A,
        16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE5D9, 16'hE5D9, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD8, 16'hDDD8, 16'hD5D8, 16'hC597, 16'hC597, 16'hC597, 16'hC598, 16'hC598, 16'hC598, 16'hC597, 16'hCDD8, 16'h93D0, 16'hA451, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hABCF, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFF1D, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9B, 16'hFE9B, 16'hF65A, 16'hDD16, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hF65B, 16'hF61A, 16'hDD16, 16'hD515, 16'hE598, 16'hF65A, 16'hF65B, 16'hEE1A, 16'hEE1A, 16'hF65A, 16'hEE1A, 16'hF65B, 16'hDD56, 16'hCC93, 16'hD4D4, 16'hDD57, 16'hF65B, 16'hEE1A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hEE1A, 16'hF65A,
        16'hCCD4, 16'hDD56, 16'hD4D4, 16'hEDD9, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hF65B, 16'hCCD4, 16'hE557, 16'hCCD4, 16'hE598, 16'hF65B, 16'hF65A, 16'hF65B, 16'hF61A, 16'hE598, 16'hD4D5, 16'hCC94, 16'hD515, 16'hEDD9, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE5D9, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD8, 16'hDDD8, 16'hD5D8, 16'hCD98, 16'hC597, 16'hC597, 16'hC597, 16'hC598, 16'hC598, 16'hC597, 16'hC598, 16'hBD15, 16'h7A8A, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD55, 16'hD596, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFEDC, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9B, 16'hF69B, 16'hF65B, 16'hFE5B,
        16'hF65A, 16'hCC94, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hF65A, 16'hE5D8, 16'hD4D4, 16'hCCD3, 16'hE597, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE1A, 16'hF65B, 16'hE598, 16'hC412, 16'hD4D4, 16'hE597, 16'hF65B, 16'hEE1A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hEE1A, 16'hF65A, 16'hD515, 16'hDD15, 16'hCC93, 16'hE598, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hF61A, 16'hF65B, 16'hDD57, 16'hE556, 16'hDD57, 16'hE597, 16'hFE5B, 16'hEDD9, 16'hD516, 16'hCC94, 16'hD4D5, 16'hE597, 16'hEE1A, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A,
        16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE5D9, 16'hE5D9, 16'hDDD9, 16'hDDD8, 16'hDDD8, 16'hDDD9, 16'hDDD9, 16'hD598, 16'hC557, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hCD98, 16'h93CF, 16'h9C50, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hABCF, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFF1D, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hF69B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF61A, 16'hD4D4, 16'hEE19, 16'hF65A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hF65A, 16'hE5D8, 16'hCC92, 16'hCC52, 16'hE598, 16'hEE1A, 16'hF65A, 16'hF65A, 16'hEE19,
        16'hC411, 16'hD493, 16'hDD57, 16'hF65B, 16'hEE1A, 16'hF65A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hEE1A, 16'hF65A, 16'hE557, 16'hD4D4, 16'hD4D5, 16'hDD56, 16'hF65B, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hF61A, 16'hF65B, 16'hF61A, 16'hDD16, 16'hE598, 16'hCC93, 16'hCC94, 16'hCC53, 16'hD4D5, 16'hEDD9, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hEE5A, 16'hF65A, 16'hE598, 16'hE5D8, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hDDD9, 16'hDDD9, 16'hDDD8, 16'hDD98, 16'hCD15, 16'hC515, 16'hC515, 16'hB493, 16'hC557,
        16'hCDD8, 16'hC598, 16'hCD98, 16'hCD98, 16'hC598, 16'hC598, 16'hBD15, 16'h7ACB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBCD3, 16'hD5D6,
        16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFEDD, 16'hFE9C, 16'hFE9B, 16'hFE5B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF61A, 16'hF61A, 16'hCCD4, 16'hEE19, 16'hF65A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hF65B, 16'hF61A, 16'hDD56, 16'hC452, 16'hC493, 16'hE557, 16'hF61A, 16'hFE5B, 16'hDD15, 16'hBBD0, 16'hDD16, 16'hF65A, 16'hEE1A, 16'hF65A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hEE1A, 16'hEE1A, 16'hF65A, 16'hEDD9, 16'hCC94, 16'hD4D5, 16'hD4D4, 16'hF65A, 16'hEE1A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF61A, 16'hE598, 16'hDCD5, 16'hC412, 16'hC452, 16'hD4D4, 16'hE597, 16'hF61A, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A,
        16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hEE1A, 16'hDD16, 16'hE5D9, 16'hF65A, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE5D9, 16'hE5D9, 16'hE619, 16'hE5D9, 16'hD557, 16'hCD15, 16'hCD56, 16'hCD15, 16'hC515, 16'hBC93, 16'hB493, 16'hB494, 16'hAC93, 16'hB4D5, 16'hA453, 16'hAC94, 16'hBD16, 16'hC557, 16'hCD98, 16'h93CF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hABCE, 16'hEE9B, 16'hF71D, 16'hEE9A, 16'hDD55, 16'hDD15, 16'hF61A, 16'hFE9C, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE1A, 16'hF61A, 16'hCCD4, 16'hE5D8, 16'hF65B, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A,
        16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hF61A, 16'hE598, 16'hCCD4, 16'hCCD4, 16'hDD16, 16'hE557, 16'hD493, 16'hDCD5, 16'hFE5B, 16'hF65B, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hF61A, 16'hF65A, 16'hEE1A, 16'hEE1A, 16'hF65A, 16'hED98, 16'hE556, 16'hD4D4, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF61A, 16'hED98, 16'hDD16, 16'hCC93, 16'hC452, 16'hD494, 16'hD4D5, 16'hEDD8, 16'hF61A, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hE597, 16'hD515, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619,
        16'hE619, 16'hE5D9, 16'hCD16, 16'hBC93, 16'hCD15, 16'hD557, 16'hCD15, 16'hBC52, 16'hA3D0, 16'hA3CF, 16'hBC93, 16'hBCD4, 16'hBCD4, 16'hC516, 16'hAC94, 16'h9C11, 16'h93D0, 16'h8B4E, 16'hACD4, 16'hAC93, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE18, 16'hAC0F, 16'hDE18, 16'hF71D, 16'hF6DC, 16'hFE5B, 16'hED98, 16'hD4D4, 16'hEDD9, 16'hFE5B, 16'hF65A, 16'hF61A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hF61A, 16'hD4D5, 16'hE598, 16'hF65B, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hF65B, 16'hF61A, 16'hEDD9, 16'hD515, 16'hD4D4, 16'hD4D4, 16'hC412, 16'hE557, 16'hEDD9, 16'hEE1A, 16'hEE5A, 16'hF65A, 16'hEE1A, 16'hEE19, 16'hF619, 16'hF619, 16'hEE19, 16'hF5D9, 16'hF5D9, 16'hDD15, 16'hE557, 16'hED98, 16'hE557, 16'hDD16, 16'hCC93, 16'hC452, 16'hC452, 16'hC452, 16'hCC94, 16'hDD56, 16'hEDD9, 16'hF65A, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A,
        16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hEE1A, 16'hD4D4, 16'hDD16, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE61A, 16'hE5D8, 16'hBC93, 16'hC494, 16'hDD97, 16'hCCD5, 16'hAC11, 16'hAC11, 16'hC4D4, 16'hD597, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hCDD8, 16'hCD98, 16'hCD98, 16'hCD98, 16'hC597, 16'hBD16, 16'h93D0, 16'h8B4E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hA3CE, 16'hBCD2, 16'hFF9E, 16'hFF9F, 16'hFEDD, 16'hFE5C, 16'hFE9C, 16'hF61A, 16'hD4D4, 16'hEDD8, 16'hF65B, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hF61A, 16'hD4D5, 16'hDD97, 16'hF65B, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A,
        16'hF65B, 16'hF65A, 16'hF65A, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hF65B, 16'hF65B, 16'hF65B, 16'hEE19, 16'hDD56, 16'hD4D4, 16'hD4D4, 16'hEE19, 16'hF65A, 16'hF65A, 16'hEE19, 16'hD4D4, 16'hB3D0, 16'hC452, 16'hC452, 16'hC411, 16'hD4D4, 16'hDCD5, 16'hD4D4, 16'hCC52, 16'hDD15, 16'hD515, 16'hDD16, 16'hE597, 16'hEE19, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hEE5A, 16'hEE1A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65B, 16'hDD57, 16'hD493, 16'hE597, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A,
        16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE619, 16'hE5D9, 16'hE619, 16'hE619, 16'hD557, 16'hBC93, 16'hD556, 16'hCD16, 16'hB411, 16'hAC10, 16'hCD15, 16'hDDD8, 16'hDDD9, 16'hD5D8, 16'hD598, 16'hD598, 16'hD598, 16'hCD98, 16'hCD98, 16'hCD97, 16'hC597, 16'hC597, 16'hCD98, 16'hCD98, 16'h9C11, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'h79C5, 16'hE659, 16'hFFDF, 16'hFF5E, 16'hF69C, 16'hF65B, 16'hF65B, 16'hFE5B, 16'hEDD9, 16'hC453, 16'hF61A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hF61B, 16'hD515, 16'hDD56, 16'hF65B, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hEDD9, 16'hEE19, 16'hEE19, 16'hEE19, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF65A, 16'hF65A, 16'hF65B,
        16'hF65B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hD4D4, 16'hD494, 16'hE5D8, 16'hF65A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hE5D9, 16'hEE1A, 16'hE5D9, 16'hC494, 16'hBC53, 16'hDD97, 16'hC493, 16'hABD0, 16'hCD15, 16'hDDD9, 16'hDDD9, 16'hD5D8, 16'hD598, 16'hD598, 16'hD598, 16'hD598, 16'hD598, 16'hCD98, 16'hCD98, 16'hCD98, 16'hCD98, 16'hCD97, 16'hC597, 16'hC597, 16'hCD97, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA410, 16'hBC92, 16'hFF5E, 16'hFFDF, 16'hFF5E, 16'hFE9C, 16'hFE5B, 16'hF65B, 16'hF61A, 16'hF65B, 16'hDD57, 16'hC452, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hF61B, 16'hD515, 16'hD515, 16'hF65B, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE5A,
        16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65B, 16'hE5D8,
        16'hCC93, 16'hD515, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hEE1A, 16'hDD97, 16'hBC11, 16'hD4D5, 16'hD557, 16'hABD0, 16'hC494, 16'hDDD9, 16'hDDD9, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD598, 16'hD598, 16'hD598, 16'hCD98, 16'hCD98, 16'hCD98, 16'hCD98, 16'hCD97, 16'hCD97, 16'hCD97, 16'hC597, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD96, 16'h8249, 16'hE659, 16'hFF9F, 16'hFFDF, 16'hFF5E, 16'hF65B, 16'hF65B, 16'hF61A, 16'hEE1A, 16'hEE1A, 16'hF61A, 16'hD515, 16'hCC93, 16'hF61A, 16'hEE1A, 16'hEE1A, 16'hEE1B, 16'hDD56, 16'hCCD4, 16'hF65B, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A,
        16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65B, 16'hD515, 16'hCC94, 16'hDD57, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hE619, 16'hEE1A, 16'hDD57, 16'hABD0, 16'hDD16, 16'hCCD4, 16'hA38F, 16'hD556, 16'hE5D9, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD598, 16'hD598, 16'hD598, 16'hCD98, 16'hCD98, 16'hCD98, 16'hCD98, 16'hCD98, 16'hCD97, 16'hC597,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hABCF, 16'hBC92, 16'hE659, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hF61A, 16'hF65A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19,
        16'hC411, 16'hE557, 16'hEE1A, 16'hEE1A, 16'hEE5B, 16'hE597, 16'hCC94, 16'hF65B, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A,
        16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE19, 16'hCCD4, 16'hCC93, 16'hDD97, 16'hF65A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hE619, 16'hEE1A, 16'hD556, 16'hC452, 16'hDD57, 16'hC453, 16'hBC52, 16'hDD98, 16'hE5D9, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hD5D8, 16'hD5D8, 16'hD598, 16'hD598, 16'hD598, 16'hD598, 16'hD598, 16'hD598, 16'hD598, 16'hCD98, 16'hCD98, 16'hCD98, 16'hCD98, 16'hCD97, 16'hCD97, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBCD2, 16'hC4D4, 16'hD556, 16'hDE59, 16'hFFDF, 16'hFF9F, 16'hFEDC, 16'hEDD9, 16'hEE19, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hE598, 16'hCC93, 16'hEDD9, 16'hEE1A, 16'hEE1A, 16'hE5D9, 16'hC453, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A,
        16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65B, 16'hDD97, 16'hCC93, 16'hD4D4, 16'hEDD9, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hE619, 16'hEE1A, 16'hDD56, 16'hC493, 16'hDD57, 16'hB411, 16'hCCD5, 16'hE5D9, 16'hDDD9, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hD5D8, 16'hD5D8, 16'hD5D8,
        16'hD598, 16'hD598, 16'hD598, 16'hD598, 16'hD598, 16'hD598, 16'hCD98, 16'hCD98, 16'hCD98, 16'hCD98, 16'hCD97, 16'hCD97, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hA34C, 16'hE619,
        16'hD556, 16'hFF9E, 16'hFF9F, 16'hFF1D, 16'hF65B, 16'hEDD9, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hD4D5, 16'hD515, 16'hF65A, 16'hEE1A, 16'hEDD9, 16'hC452, 16'hEE19, 16'hEE5A, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A,
        16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hD514, 16'hD514, 16'hD4D4, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE619, 16'hEE1A, 16'hDD56, 16'hBC52, 16'hDD16, 16'hBC12, 16'hD516, 16'hE61A, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD598, 16'hD598, 16'hD598, 16'hD598, 16'hD598, 16'hD598, 16'hCD98, 16'hCD98, 16'hCD98, 16'hCD98, 16'hCD98, 16'hCD97, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBC91, 16'hD556, 16'hE619, 16'hD556, 16'hFF9E, 16'hFF1C, 16'hFE9C, 16'hF61A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEDD9, 16'hBC11, 16'hDD97, 16'hEE5B, 16'hEE1A, 16'hC452, 16'hE5D9, 16'hF65A, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B,
        16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hEE19, 16'hCC93, 16'hD514, 16'hCCD4, 16'hF65B, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE19, 16'hEE1A, 16'hDD56, 16'hC452, 16'hD516, 16'hC493, 16'hDD98,
        16'hE61A, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD598, 16'hD598, 16'hD598, 16'hCD98, 16'hCD98, 16'hCD98, 16'hCD98, 16'hCD98, 16'hCD98, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'h9B0B, 16'hF6DB, 16'hD556, 16'hF69B, 16'hFF1D, 16'hFEDC, 16'hFE9C, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE1A, 16'hDD56, 16'hCC94, 16'hEE1A, 16'hF61B, 16'hCC93, 16'hE598, 16'hF65B, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF61A, 16'hEE1A, 16'hF65A, 16'hF65A, 16'hF65A,
        16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65B, 16'hDD56, 16'hD4D4, 16'hCCD4, 16'hE598, 16'hF65B, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hDD97, 16'hBC53, 16'hD516, 16'hC4D4, 16'hE5D9, 16'hE5DA, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hD598, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD598, 16'hD598, 16'hD598, 16'hCD98, 16'hCD98, 16'hCD98, 16'hCD98, 16'hCD98, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC514, 16'hDDD7, 16'hFF1D, 16'hBBD1, 16'hF69B, 16'hFE9B, 16'hFE9B, 16'hF65A, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hEE19, 16'hF61A, 16'hC493, 16'hDD57, 16'hF65B, 16'hCC94, 16'hDD56, 16'hF65B, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A,
        16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65B, 16'hDD15, 16'hE597, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5B, 16'hF65A, 16'hF65A, 16'hF65A, 16'hF65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hF65B, 16'hCCD3, 16'hDD15, 16'hCC93, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE1A,
        16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hE5D8, 16'hC493, 16'hD557, 16'hD556, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD598, 16'hD598, 16'hCD98, 16'hCD98, 16'hCD98, 16'hCD98, 16'hCD98
    };

    reg [15:0] image_succeeded [0:65535] = {
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hAD55, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h8410, 16'h7BCF, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h8C51, 16'h8C51, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hAD55, 16'hBDD7, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8C51, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8410, 16'h7BCF, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8410, 16'h9492, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h9492, 16'h9492, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8C51, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h8410, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8410, 16'h9492, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hDEDB, 16'hD69A, 16'hD69A, 16'hD69A, 16'hE71C, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hB596, 16'h9492, 16'h8410, 16'h8410, 16'h8410, 16'h8410, 16'h8C51, 16'h9492, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h8C51, 16'h9492, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51,
        16'h9492, 16'h8410, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h8410, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8C51, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hEF5D, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h8C51, 16'h9492, 16'h9492, 16'h8410, 16'h8C51, 16'h8C51, 16'h8410, 16'h8410, 16'h8410, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8410, 16'h9492, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h8C51, 16'h9492, 16'h9CD3, 16'hBDD7, 16'hAD55, 16'h9CD3, 16'h8C51, 16'h8410, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h8C51, 16'h9CD3, 16'hCE59, 16'hE71C, 16'hEF5D, 16'hDEDB, 16'hCE59, 16'hBDD7, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'hC618, 16'hAD55, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8451, 16'h9492, 16'h8C51, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h8410,
        16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hEF5D, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h7BCF, 16'h8C51, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'h8C51, 16'h7BCF, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8C51, 16'h9492, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h9492, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hC618, 16'hA514, 16'h9492, 16'h9492, 16'h8C51, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h8C51, 16'h9CD3, 16'h9492, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h9CD3, 16'hB596, 16'hC618, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8C51, 16'h9492, 16'h8C51, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8C51, 16'h9492, 16'h9CD3, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hBDD7, 16'h8C51, 16'h8410, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h8410, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8C51, 16'h8C51, 16'h9CD3, 16'hA514, 16'h9492, 16'h9492, 16'h8C51, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8410, 16'h9492, 16'h8C51, 16'h9492, 16'hC618, 16'hDEDB, 16'hE71C, 16'hEF5D, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8C51, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'hB596, 16'hA514, 16'hA514, 16'hB596, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hA4D3, 16'h8410, 16'h9492, 16'h9CD3, 16'h9492, 16'h8C51, 16'h9492, 16'h9492, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hEF5D, 16'hFFDF, 16'hF79E, 16'h9CD3, 16'h9492, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h8C51, 16'h9492, 16'h9492, 16'h8410, 16'h8410, 16'h8C51, 16'h9492, 16'h9CD3, 16'hAD55, 16'hC618, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h7BCF, 16'h8C51, 16'h8C51, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hB596, 16'h8410, 16'h8C51, 16'h9492, 16'h8C51, 16'h8C51, 16'h8410, 16'hA514, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9CD3, 16'h8C51, 16'h9492, 16'h9492, 16'h8410, 16'h9CD3, 16'hAD55, 16'h9492, 16'h9492, 16'h8410, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8C51, 16'h9492, 16'h9CD3, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h9492, 16'h8410, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'h8410, 16'h8C51, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'hA514, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hA514, 16'h8410, 16'h9492, 16'h9492, 16'h8C51, 16'h8C51, 16'h9492, 16'h9CD3, 16'h8410, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'hC618, 16'hF79E, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8410, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hC618, 16'h9CD3, 16'h8C51, 16'h8410, 16'h8410, 16'h8410, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h8410, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8C51, 16'h8C51, 16'h9CD3, 16'hCE59, 16'hA514, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'hAD55, 16'hAD55, 16'h8C51, 16'h8C51, 16'h8410, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8410, 16'h9492, 16'h9492, 16'h9492, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h8C51, 16'h8C51, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h9492, 16'h8410, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hDEDB, 16'hD69A, 16'hC618, 16'hAD55, 16'h8C51, 16'h8C51, 16'h9492, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h8C51, 16'h9492, 16'h8C51, 16'h8410, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hAD55, 16'hA514, 16'hEF5D, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'hE71C,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8C51, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h8410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h9CD3, 16'h8C51, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hCE59, 16'hBDD7, 16'hBDD7, 16'hD69A, 16'hEF5D, 16'hFFDF, 16'hE71C, 16'hA514, 16'hAD55, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8410, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h9492, 16'h8410, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8410, 16'h9492, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h9492, 16'h8410, 16'hDEDB,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8C51, 16'h9492, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hAD55, 16'h8C51, 16'h8410, 16'h8C51, 16'h8410, 16'h8410, 16'h8C51, 16'hB596, 16'h9CD3, 16'h8C51, 16'h8410, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h9CD3, 16'h9492, 16'h9492, 16'h9492, 16'h8410, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8C51, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h9CD3, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h8C51, 16'h8C51, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h7BCF, 16'h9492, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hEF5D, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h8C51, 16'h9492, 16'h9CD3, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8C51, 16'h9492, 16'h8C51, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8C51, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h7BCF, 16'h8410,
        16'hAD55, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8C51, 16'h9492, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hBDD7, 16'h9CD3, 16'h9492, 16'h9492, 16'hB596, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'hB596, 16'h9CD3, 16'h9492, 16'h9492, 16'hA514, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h9492, 16'h8C51, 16'h8410, 16'h8C51, 16'h9492, 16'h8410, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8410, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h8410, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9CD3, 16'h9492, 16'h8C51, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8410, 16'h9492, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h8C51, 16'h9492, 16'h8C51, 16'h8C51, 16'hB596, 16'hD69A, 16'hE71C, 16'hE71C, 16'hB596, 16'h8C51, 16'h9492, 16'h8C51, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8410, 16'h8C51, 16'h8410, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hBDD7, 16'h8C51, 16'h8410, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'h8C51, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hAD55, 16'h8410, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'h8410, 16'hA514, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'h9D14, 16'hD69A, 16'hEF5D, 16'hEF5D, 16'hDEDB, 16'hB596, 16'h8C51, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h9492, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8C51, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492,
        16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h7BCF, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'h8410, 16'h8C51, 16'h8410, 16'h8C51, 16'h9492, 16'h9492, 16'h8410, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hB596, 16'hBDD7, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h9492, 16'h8410, 16'h9492, 16'h9492, 16'h9492, 16'h8410, 16'h9492, 16'h9492, 16'h9492, 16'h8410, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h8410, 16'hC618, 16'hE71C, 16'h9492, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'h8C51, 16'h9492, 16'h9492, 16'h8410, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8410, 16'h9492, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hAD55, 16'h8C51, 16'h9492, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h8410, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h9492, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h9492, 16'h8410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h8410, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8C51, 16'h8410, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h8410, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8410, 16'h9492, 16'h9492, 16'h9492, 16'h8410, 16'h9CD3, 16'hBDD7, 16'h9CD3, 16'h8C51,
        16'h9CD3, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8410, 16'h9492, 16'h8C51, 16'h8C51, 16'h8C51, 16'h9492, 16'h9492, 16'h8410, 16'h9CD3, 16'hBDD7, 16'hBDD7, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h8410, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492,
        16'h8C51, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9CD3, 16'h9492, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hC618, 16'h9CD3, 16'h8C51, 16'h8410, 16'h8410, 16'h8410, 16'h8410, 16'h9492, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hAD55, 16'h8410, 16'h9492, 16'h9492, 16'h8C51, 16'h9492, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9CD3, 16'h8410, 16'h8410, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hC618, 16'hAD55, 16'h9CD3, 16'h9CD3, 16'hB596, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8410, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'h9492, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8410, 16'h9492, 16'h8410, 16'hD69A,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h8410, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h9492, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h8C51, 16'h9492, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h8410, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8C51, 16'h9492, 16'h9CD3, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hDEDB, 16'hD69A, 16'hD69A, 16'hDEDB, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hA514, 16'h8C51, 16'h9492, 16'h9492, 16'h8410, 16'hAD55, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hB596, 16'hAD55, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8C51, 16'h8410, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'h8410, 16'hAD55, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8410, 16'h9492, 16'h8410, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8C51, 16'h9492, 16'h9CD3, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8C51, 16'h9492, 16'h9492, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492,
        16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h8410, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8410, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDE, 16'hF75E, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8410, 16'h9492, 16'h9492, 16'h8410, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8410, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'h9CD3, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h9492, 16'h9492,
        16'h8410, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8410, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8410, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8410, 16'h9492, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8410, 16'h9492, 16'h8C51, 16'hA514, 16'hE71C, 16'hF79E, 16'hF79E, 16'hE71C, 16'hC618, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h9CD3, 16'h8C51, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hC596, 16'h93CF, 16'h7B0C, 16'h7B0C, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h9492, 16'h9492, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8410, 16'h9492, 16'h9492, 16'h8410, 16'h9492, 16'hAD55, 16'h9D14, 16'h8410, 16'h9492, 16'h9492, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h8C51, 16'h9492, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h8C51, 16'h9492, 16'h9CD3, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8410, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h9492, 16'h8410, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h8410,
        16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'h8410, 16'h9492, 16'h9492, 16'h8C51, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'hAD55, 16'hAD55, 16'h8410, 16'h9492, 16'h8410, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hDE9A, 16'hA492, 16'h51C6, 16'h3000, 16'h2800, 16'h800, 16'h000, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h9451, 16'h9492, 16'h8410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h9492, 16'h9492, 16'h8C51, 16'hC618, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8C51,
        16'h9492, 16'h9492, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8C51, 16'h9492, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8C51, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h9CD3, 16'h8410, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h8410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h8410, 16'h9CD3, 16'hF79E, 16'hFFDF, 16'hB596, 16'h9492, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hDE9B, 16'hBD55, 16'h834D, 16'h7A8B, 16'h5946, 16'h4104, 16'h4986, 16'h5186, 16'h5A08, 16'h000, 16'hC5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h9492, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9CD3, 16'h9492, 16'h9492, 16'h8C51, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8C51, 16'h9492, 16'h8C51, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8410, 16'h9492, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8410, 16'h9492, 16'h8410, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492,
        16'h9492, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h9492, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h9CD3, 16'h8410, 16'h8C51, 16'h8C51, 16'h8410, 16'h8410, 16'h8C51, 16'h9492, 16'hBDD7, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'hBD96, 16'h7B0D, 16'h6A0A, 16'h830D, 16'hA452, 16'h8B8F, 16'h51C7, 16'h8B0B, 16'h9B4C, 16'hABCE, 16'hB410, 16'h5800, 16'hC5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8C51, 16'h9492, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hD69A, 16'h8410, 16'h9492, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8C51, 16'h9492, 16'h8410, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h9492, 16'h8410, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h8410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h9492, 16'h9492, 16'h9492, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8C51, 16'h9492, 16'h9CD3, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hD69A, 16'hBDD7, 16'hB596, 16'hC618, 16'hD69A, 16'hE71C, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hC596, 16'h7B4C, 16'h59C8, 16'h830E, 16'hA452, 16'hB4D4, 16'hC556, 16'hA452, 16'h5185, 16'hAB8E, 16'hC451, 16'hC451, 16'hC451, 16'hCC92, 16'h79C7, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8C51, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8410, 16'h9492, 16'h8410, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h8410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h8410, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8410, 16'h9492,
        16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hA514, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8C51, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hC596, 16'h8B8E, 16'h6208, 16'h6A4B, 16'h93D0, 16'hAC94, 16'hBD15, 16'hBCD5, 16'hC516, 16'hA452, 16'h51C7, 16'hABCF, 16'hCC51, 16'hC451, 16'hC451, 16'hBC51, 16'hC492, 16'h8208, 16'hB555, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h8410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9CD3, 16'h9492, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h9CD3, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h7BCF, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hBD96, 16'h9C51, 16'h8B4D, 16'h7ACC, 16'h9390, 16'hAC93, 16'hBD15, 16'hBD16, 16'hBD15, 16'hB4D4, 16'hBD16, 16'h9C11, 16'h5986, 16'hAC0F, 16'hC452, 16'hC451, 16'hC451, 16'hC451, 16'hC451,
        16'hCC92, 16'h8208, 16'hBD56, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h9492, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h8410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h9492, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h8C51, 16'h8C51, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hAD55, 16'h8C51, 16'h9492, 16'h9CD3, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8410, 16'h9492, 16'h9492, 16'h8C51, 16'hA514, 16'hBDD7, 16'hC618, 16'hBDD7, 16'h9CD3, 16'h8410, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h9492, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hBD56, 16'h9BCF, 16'h9B8F, 16'hB514, 16'hD659, 16'hCD96, 16'hC515, 16'hBD15, 16'hBD15, 16'hB4D5, 16'hBCD5, 16'hB4D5, 16'hBD15, 16'h9C52, 16'h61C8, 16'hB40F, 16'hCC91, 16'hC451, 16'hC451, 16'hC451, 16'hBC51, 16'hC451, 16'hCC92, 16'h8A49, 16'hB555, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hCE59, 16'h8410, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h9492, 16'h8410, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h9492, 16'h8C51, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8C51, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8410, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8410, 16'h9492, 16'h9492, 16'h8C51, 16'h8C51, 16'h8410, 16'h8C51, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'h8C51, 16'h9492, 16'h9492, 16'h8410, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hBD96, 16'h9C10, 16'h938E, 16'hBD56, 16'hEEDC, 16'hF75D, 16'hEEDC, 16'hC556, 16'hB4D4, 16'hBD15, 16'hBCD5, 16'hBD15, 16'hBD15,
        16'hBCD5, 16'hBD15, 16'hAC53, 16'h59C7, 16'hB410, 16'hC491, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hCC92, 16'h8A49, 16'hB514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8410, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h8C51, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h9492, 16'h9492, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hCE59, 16'h8410, 16'h9492, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h9492, 16'h8410, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8410, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'h8410, 16'h8410, 16'hB596, 16'hE71C, 16'h9CD3, 16'h9492, 16'h8C51, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hC596, 16'h8B4D, 16'h8B8E, 16'hB4D4, 16'hE69A, 16'hFF9E, 16'hFF5E, 16'hDE5A, 16'hBD15, 16'hB494, 16'hBCD4, 16'hBD15, 16'hBD15, 16'hBCD5, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBCD5, 16'h6209, 16'hABCF, 16'hCC92, 16'hC451, 16'hC491, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hCC92, 16'h8A49, 16'hBD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8410, 16'h9492, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h8410, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h8410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h8410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'hAD55, 16'h9492, 16'h8C51, 16'h8C51, 16'h9492, 16'hA514, 16'hC618, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h8C51, 16'h8C51, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hCE18, 16'h93CF, 16'h7A8A, 16'hB4D3, 16'hE6DB, 16'hFF9F, 16'hFF9F,
        16'hEEDC, 16'hCD98, 16'hB4D4, 16'hB494, 16'hBCD5, 16'hC516, 16'hBD16, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBCD5, 16'hBD15, 16'h7B0D, 16'h934D, 16'hCC92, 16'hC451, 16'hC491, 16'hC491, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hCC92, 16'h8208, 16'hBD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h8410, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8C51, 16'h9492, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h8410, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hEF5D, 16'hEF5D, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8C51, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h9C10, 16'h824B, 16'h938F, 16'hD658, 16'hFF9E, 16'hFFDF, 16'hF71D, 16'hD619, 16'hBD15, 16'hB493, 16'hB4D5, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD16, 16'hBD15, 16'hBD15, 16'hBD16, 16'hC556, 16'h93D0, 16'h7A8A, 16'hC492, 16'hC451, 16'hC491, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC492, 16'hD514, 16'h8249, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h9492, 16'h9492, 16'h8C51, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hB596, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9CD3, 16'h9492, 16'h9492, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h8C51, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9CD3, 16'h9492, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h7BCF, 16'h8410, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8410, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFF9E, 16'hF79E, 16'hF79D, 16'hF79E, 16'hF79E, 16'hFF9E, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB,
        16'hB514, 16'h934E, 16'h93CE, 16'hCD97, 16'hF75D, 16'hFFDF, 16'hFF9E, 16'hE69A, 16'hC516, 16'hB494, 16'hB4D5, 16'hBD15, 16'hBD16, 16'hBD16, 16'hBD16, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hC516, 16'hBD15, 16'hBD16, 16'hC556, 16'hA452, 16'h7249, 16'hBC51, 16'hC491, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC492, 16'hD4D4, 16'hDD55, 16'h8A4A, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h8C51, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h7BCF, 16'h9492,
        16'h8410, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8C51, 16'h9492, 16'h8C51, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9CD3, 16'h8C51, 16'h9492, 16'h8410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8C51, 16'h8C51, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hEF1C, 16'hD659, 16'hCD97, 16'hCD96, 16'hBCD4, 16'hA410, 16'hAC92, 16'hCD97, 16'hD597, 16'hD5D8, 16'hA411, 16'h834D, 16'h7B0C, 16'h72CB, 16'h6A8A, 16'h72CA, 16'h72CB, 16'h7B0C, 16'h7B0C, 16'h8B8E, 16'h93CF, 16'hA492, 16'hAD14, 16'hC5D7, 16'hD699, 16'hE6DB, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hC596, 16'h8B4D, 16'h8B4D, 16'hBD55, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hD598, 16'hBCD5, 16'hB4D5, 16'hBD16, 16'hBD16, 16'hC556, 16'hBD16, 16'hBD16, 16'hBD16, 16'hBD16, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hC516, 16'hB493, 16'h724A, 16'hB410, 16'hC492, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hCCD3, 16'hD514, 16'hDD55, 16'h8A4A, 16'hC596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8410, 16'h9492, 16'h8410, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'hC618, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h9CD3, 16'h8C51, 16'h9492, 16'h8C51, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8C51, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hD659, 16'hC556, 16'hBD14, 16'hAC92, 16'hB492, 16'hAC52, 16'hB4D3, 16'hCDD7, 16'hDE59, 16'hE69B, 16'hEF1C, 16'hEEDC, 16'hDE5A, 16'hCD56, 16'hAC52, 16'h9BD0, 16'hA452, 16'hA452, 16'hB493, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB494, 16'hAC93, 16'hAC53, 16'h9C11, 16'h9390, 16'h8B8F, 16'h72CB, 16'h6A49, 16'h61C7, 16'h6A4A, 16'h7B4D, 16'h9C51, 16'hC596, 16'hDE9B, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE5A, 16'hA411, 16'h7A8A, 16'hAC92, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hDE19, 16'hC515, 16'hBCD5, 16'hBD15, 16'hBD16, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hBD16, 16'hBD16, 16'hC516, 16'hBD16, 16'hBD16, 16'hBD16, 16'hBD15, 16'hBD16, 16'hBD15, 16'hC516, 16'hBCD4, 16'h7249, 16'hABCF, 16'hCC92, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hCC93, 16'hDD14, 16'hDD15, 16'hDD55, 16'h8208, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'hDEDB, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8410, 16'h9492, 16'h8410, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8410, 16'h9492, 16'h9492, 16'h8410, 16'h9492, 16'hAD55, 16'hA514, 16'h8C51, 16'h8C51, 16'h9492, 16'h9492, 16'h8410, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8C51, 16'h9492, 16'h8C51, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hD618, 16'hB4D3, 16'hA3D0, 16'hA410, 16'hBD14, 16'hCDD8, 16'hE6DB, 16'hF75D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hE69A, 16'hBD14, 16'hAC52, 16'hAC93, 16'hBCD5, 16'hBCD4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB514, 16'hB514, 16'hB4D4, 16'hBD15, 16'hBD56, 16'hC556, 16'hCD97, 16'hC556, 16'hCD97, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hC597, 16'hB515, 16'h9411, 16'h7B0C, 16'h6208, 16'h59C7, 16'h7B4D, 16'hAD14, 16'hDE9A, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hC556, 16'h828B, 16'h7249, 16'hBD55, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'hCD97, 16'hBCD5, 16'hBCD5, 16'hBD15, 16'hC516, 16'hC516, 16'hC556, 16'hC556, 16'hBD16, 16'hBD16, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC516, 16'hBD15, 16'hBD15, 16'hC516, 16'hC516, 16'h8B4E, 16'hA38E, 16'hC492, 16'hC451, 16'hC492, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451,
        16'hCC92, 16'hDD14, 16'hDD15, 16'hDD15, 16'hDD15, 16'h79C7, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8410, 16'h9492, 16'h9492, 16'h9492, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8410, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'hBDD7, 16'hDEDB, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hBDD7, 16'h8C51, 16'h9492, 16'h9492, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hDE5A, 16'hB4D3, 16'h938E, 16'hA3CF, 16'hBCD3, 16'hDE59, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hD598, 16'hBD15, 16'h9BD0, 16'hAC52, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hBCD4, 16'hBCD4, 16'hBD14, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hBD14, 16'hBD15, 16'hC556, 16'hC556, 16'hC556, 16'hCD97, 16'hD619, 16'hDE19, 16'hDE1A, 16'hDE5A,
        16'hDE5A, 16'hDE5A, 16'hDE19, 16'hCD97, 16'hAC93, 16'h830D, 16'h4904, 16'h628A, 16'hA492, 16'hDE9A, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hD618, 16'hA451, 16'h6186, 16'h938D, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hDE19, 16'hCD56, 16'hBCD5, 16'hBD15, 16'hBD56, 16'hC556, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hC556, 16'hC516, 16'hC516, 16'hC556, 16'hBD56, 16'hC556, 16'hC556, 16'hC516, 16'hC516, 16'hBD16, 16'hBD16, 16'hC516, 16'hC516, 16'h938F, 16'hB451, 16'hC492, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hD4D4, 16'hDD15, 16'hDD15, 16'hDD15, 16'hDD15, 16'h7186, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'hC618, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hC618, 16'h8C51, 16'h9492, 16'h9492, 16'h8410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8C51, 16'h8410, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'h8410, 16'h9CD3, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h7BCF, 16'h8C51, 16'h8410, 16'h9492, 16'hAD55, 16'hBDD7, 16'hB596, 16'hA514, 16'h8C51, 16'h8C51, 16'h9492, 16'h9492, 16'h8410, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE5A, 16'hB4D3, 16'h938E, 16'hA410, 16'hCD96, 16'hEEDB, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF75D, 16'hF6DD, 16'hEE9B, 16'hE65A, 16'hEE9C, 16'hE65A, 16'hBCD4, 16'hA411, 16'h938F, 16'hA3D0, 16'hAC52, 16'hB452, 16'hAC53, 16'hAC93, 16'hB4D4, 16'hBD15, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hCD97, 16'hD5D8, 16'hDE19, 16'hDE19, 16'hDE1A, 16'hDE19, 16'hDE5A, 16'hDE5A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hD619, 16'hBD15, 16'h8B4E, 16'h61C7, 16'h72CB, 16'hAC93, 16'h9B8F, 16'h9BCF, 16'hD5D7, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hF6DC, 16'hD597, 16'hC4D5, 16'hBCD5, 16'hC516, 16'hC556, 16'hBD16, 16'hC516, 16'hC556, 16'hC516, 16'hC516, 16'hC516, 16'hC556, 16'hC556, 16'hC516, 16'hC516, 16'hC556, 16'hBD16, 16'hC516, 16'hC516, 16'hC556, 16'hBD16, 16'hC516, 16'hC516, 16'hC556, 16'h9BD0,
        16'h9C51, 16'hD5D7, 16'hC514, 16'hC492, 16'hC451, 16'hC491, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hD4D3, 16'hDD15, 16'hDD15, 16'hDD15, 16'hDD15, 16'hDD14, 16'h7187, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9CD3, 16'h8C51, 16'h9492, 16'h9492, 16'h8410, 16'h9492, 16'hAD55, 16'hBDD7, 16'hB596, 16'h9492, 16'h8410, 16'h9492, 16'h9492, 16'h8410, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hBDD7, 16'hA514, 16'h9CD3, 16'h9CD3, 16'hAD55, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8410, 16'h9CD3, 16'h9492, 16'h9492, 16'h8C51, 16'h8C51, 16'h8C51, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h8410, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hC555, 16'h9B8E, 16'hA3CF, 16'hCD96, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hF6DB, 16'hCD15, 16'hAC12, 16'hB452, 16'hB493, 16'hBC94, 16'hC516, 16'hB493, 16'hAC52, 16'hBCD4, 16'hBD15, 16'hC515, 16'hB4D4, 16'hA411, 16'h9BCF, 16'h9B8F, 16'hB493, 16'hD5D8, 16'hE65A, 16'hDE5A,
        16'hDE5A, 16'hDE5A, 16'hDE1A, 16'hDE19, 16'hD619, 16'hCDD8, 16'hCD98, 16'hCD97, 16'hCDD8, 16'hD5D8, 16'hDE19, 16'hDE5A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE5A, 16'hDE19, 16'hDE19, 16'hDE5A, 16'hE69B, 16'hEE5A, 16'h934D, 16'h4800, 16'hB514, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFF5D, 16'hE65A, 16'hD557, 16'hC515, 16'hBD15, 16'hC516, 16'hBD16, 16'hC556, 16'hC556, 16'hBD16, 16'hC556, 16'hC556, 16'hC516, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hBD16, 16'hC557, 16'hA452, 16'h8BCF, 16'hCE17, 16'hC617, 16'hD658, 16'hD5D7, 16'hC514, 16'hC451, 16'hC451, 16'hC452, 16'hC451, 16'hC451, 16'hCCD3, 16'hDD14, 16'hDD15, 16'hDD15, 16'hDD15, 16'hDD15, 16'hD4D4, 16'h7249, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h9CD3, 16'h8410, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'h8C51, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h8410, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hAD55, 16'h8C51, 16'h8410, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'h8C51, 16'h8410, 16'h9492, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE5A, 16'hA451, 16'h92CC, 16'hBD55, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5E, 16'hDE19, 16'hB493, 16'hAC52, 16'hBCD4, 16'hBCD4, 16'hB493, 16'hB493, 16'hC515, 16'hDDD8, 16'hDE19, 16'hDE1A, 16'hDE5A, 16'hDE19, 16'hCD97, 16'hC556, 16'hB493, 16'hA3D0, 16'h934D, 16'h934E, 16'hB493, 16'hD5D8, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65B, 16'hE65B, 16'hE65A, 16'hDE59, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE5A, 16'hDE5A, 16'hE65A, 16'hE65A, 16'hDE5A, 16'hDE5A, 16'hD619, 16'hCD56, 16'h8B0D, 16'hB4D3, 16'hFF5D, 16'hFFDF, 16'hFF9E, 16'hEE9A, 16'hD556, 16'hCCD4, 16'hBCD4, 16'hBCD5, 16'hC516, 16'hC516, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC516, 16'hC556, 16'hC516, 16'hC556,
        16'hC556, 16'hC556, 16'hC516, 16'hBD16, 16'hC516, 16'hC516, 16'hC516, 16'hC515, 16'hC556, 16'hAC93, 16'h8B8F, 16'hC5D7, 16'hC658, 16'hCE98, 16'hD69A, 16'hD69A, 16'hD659, 16'hCD96, 16'hC451, 16'hC451, 16'hC492, 16'hCC92, 16'hDD14, 16'hDD55, 16'hDD15, 16'hDD15, 16'hDD15, 16'hE556, 16'hC452, 16'h72CB, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h9492, 16'h8410, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'h8410, 16'h8C51, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hCE59, 16'hAD55, 16'h9CD3, 16'h9492, 16'h9CD3, 16'hA514, 16'hB596, 16'hD69A, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD618, 16'h9B8F, 16'h9B4E, 16'hD5D7, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hEE9C, 16'hDE19, 16'hDDD9, 16'hE61A, 16'hDDD9, 16'hBC93, 16'hAC52, 16'hBCD4, 16'hBD15, 16'hBCD4, 16'hB4D4, 16'hBCD4, 16'hB493, 16'hB4D4, 16'hD5D8,
        16'hD619, 16'hDE19, 16'hDE1A, 16'hDE19, 16'hCD97, 16'hCD97, 16'hCD97, 16'hC556, 16'hBD15, 16'hAC52, 16'h9BCF, 16'h9BD0, 16'hC556, 16'hDE5A, 16'hE65A, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE5A, 16'hDE5A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE19, 16'hB452, 16'hCD97, 16'hFFDF, 16'hEEDC, 16'hD597, 16'hC4D5, 16'hC4D5, 16'hC515, 16'hBD15, 16'hC516, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hC556, 16'hB4D4, 16'h834E, 16'hC5D7, 16'hC658, 16'hD699, 16'hDEDA, 16'hD69A, 16'hD699, 16'hD699, 16'hD69A, 16'hD5D7, 16'hC492, 16'hCC92, 16'hD514, 16'hDD15, 16'hDD15, 16'hDD15, 16'hDD15, 16'hDD15, 16'hE556, 16'hB411, 16'h834D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hCE59, 16'hAD55, 16'h9CD3, 16'h9CD3, 16'hA514, 16'hAD55, 16'hC618, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hF79E, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCDD8, 16'h930D, 16'hA3CF, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hF71D, 16'hDE19, 16'hCD56, 16'hC515, 16'hC556, 16'hC516, 16'hBC94, 16'hB493, 16'hBCD4, 16'hBD15, 16'hBCD4, 16'hB493, 16'hB494, 16'hBCD4, 16'hBCD4, 16'hAC53, 16'hBCD4, 16'hCD97, 16'hCD97, 16'hDE19, 16'hDE1A, 16'hDE1A, 16'hDE1A, 16'hCD97, 16'hC556, 16'hC597, 16'hCD97, 16'hCD57, 16'hC556, 16'hB4D4, 16'hA411, 16'hBD15, 16'hCD98, 16'hD598, 16'hDE1A, 16'hE65B, 16'hE69B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDDD9, 16'hCD57, 16'hC516, 16'hBCD4, 16'hBCD4, 16'hBD15, 16'hBD15, 16'hC515, 16'hC516, 16'hC516, 16'hC556, 16'hC556, 16'hC556,
        16'hCD57, 16'hCD57, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC516, 16'hC516, 16'hC556, 16'hBCD5, 16'h834D, 16'hBD96, 16'hCE99, 16'hD69A, 16'hE6DB, 16'hDEDB, 16'hDE9A, 16'hD699, 16'hD699, 16'hD69A, 16'hDE9A, 16'hD618, 16'hD555, 16'hDD15, 16'hDD15, 16'hDD15, 16'hDD15, 16'hDD15, 16'hDD15, 16'hE556, 16'hA34E, 16'h9C51, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD618, 16'h8ACC, 16'hA3D0, 16'hE69B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hF6DC, 16'hFF9E, 16'hFFDF, 16'hF6DD, 16'hD557, 16'hB494, 16'hBCD4, 16'hC556, 16'hCD56, 16'hC515, 16'hBCD4,
        16'hC515, 16'hC516, 16'hC515, 16'hBCD4, 16'hB493, 16'hC515, 16'hC556, 16'hBCD4, 16'hBD15, 16'hB493, 16'hBD15, 16'hD598, 16'hC557, 16'hD5D8, 16'hDE1A, 16'hDE1A, 16'hE65A, 16'hDE19, 16'hCD97, 16'hCD57, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hC557, 16'hBD15, 16'hD5D8, 16'hC556, 16'hBCD5, 16'hCD57, 16'hDE19, 16'hE65A, 16'hE69B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE69B, 16'hE69B, 16'hE65A, 16'hE65B, 16'hDE19, 16'hC556, 16'hBD16, 16'hC516, 16'hC556, 16'hC515, 16'hC515, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC557, 16'hCD57, 16'hCD57, 16'hC556, 16'hC556, 16'hC556, 16'hC557, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC516, 16'hC516, 16'hBD15, 16'h8B8F, 16'hBD96, 16'hD699, 16'hD699, 16'hD69A, 16'hDEDB, 16'hDEDB, 16'hDEDA, 16'hDE9A, 16'hCE17, 16'hC596, 16'hCDD7, 16'hD5D7, 16'hD596, 16'hD514, 16'hDD15, 16'hDD15, 16'hDD15, 16'hDD15, 16'hDD15, 16'hE556, 16'h9B0D, 16'h9C91, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69B, 16'hA38F, 16'h92CC, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF1D, 16'hEE9B, 16'hF69C, 16'hFF5E, 16'hFF5E, 16'hDE19, 16'hBC93, 16'hBCD4, 16'hC516, 16'hCD56, 16'hCD56, 16'hCD56, 16'hBCD4, 16'hC516, 16'hCD56, 16'hC515, 16'hC515, 16'hB494, 16'hC515, 16'hDE1A, 16'hD5D8, 16'hBD15, 16'hC515, 16'hB493, 16'hC516, 16'hD5D8, 16'hCD97, 16'hCD97, 16'hDE19, 16'hDE1A, 16'hDE1A, 16'hE65A, 16'hD619, 16'hCD98, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD98, 16'hD5D8, 16'hD5D8, 16'hE65A, 16'hC556, 16'hB4D4, 16'hBCD5, 16'hCD56, 16'hDE19, 16'hE65B, 16'hE65A, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65A, 16'hE69B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A,
        16'hE69B, 16'hE65A, 16'hCD97, 16'hBCD4, 16'hBCD5, 16'hC515, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hCD57, 16'hCD57, 16'hCD97, 16'hCD57, 16'hCD57, 16'hC557, 16'hC556, 16'hC557, 16'hC557, 16'hC556, 16'hC556, 16'hC557, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC516, 16'h938F, 16'hB595, 16'hD69A, 16'hD699, 16'hCE59, 16'hE71C, 16'hEF1C, 16'hDE9A, 16'hDEDA, 16'hDEDA, 16'hD658, 16'hBC92, 16'hC492, 16'hC492, 16'hCC93, 16'hD514, 16'hDD55, 16'hDD55, 16'hDD55, 16'hDD15, 16'hDD15, 16'hE556, 16'h8209, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFF9E, 16'hF75D, 16'hEF1D, 16'hF75E, 16'hF75D, 16'hEF5D, 16'hEF1C, 16'hEF1C, 16'hEF1C, 16'hEF1D, 16'hEF5D, 16'hF75D, 16'hF75D, 16'hF75E, 16'hF79E, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFF9E, 16'hEF5D, 16'hEF1C, 16'hE6DB, 16'hDE9A, 16'hDE59, 16'hBD55, 16'hC596, 16'hA411, 16'h7208, 16'hC596, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hEE9B, 16'hE65A, 16'hF69C,
        16'hFF1D, 16'hE65A, 16'hBCD4, 16'hB493, 16'hBD15, 16'hCD56, 16'hC556, 16'hCD56, 16'hCD97, 16'hC515, 16'hC556, 16'hCD97, 16'hCD56, 16'hC556, 16'hBD15, 16'hC515, 16'hE65A, 16'hE65B, 16'hDE19, 16'hC556, 16'hC515, 16'hBCD4, 16'hCD97, 16'hD5D8, 16'hCD97, 16'hCD97, 16'hD5D9, 16'hDE1A, 16'hDE1A, 16'hDE5A, 16'hE65A, 16'hDE19, 16'hCD97, 16'hCD97, 16'hCD98, 16'hCD98, 16'hD5D8, 16'hD619, 16'hD5D9, 16'hDE1A, 16'hE65A, 16'hCD97, 16'hBD15, 16'hBD15, 16'hBD15, 16'hD5D8, 16'hEE9B, 16'hE65A, 16'hDE1A, 16'hE69B, 16'hE65B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hDDD8, 16'hC515, 16'hB493, 16'hBD15, 16'hC556, 16'hC556, 16'hCD97, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD57, 16'hC557, 16'hC557, 16'hC557, 16'hC556, 16'hC516, 16'hC556, 16'hC557, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hCD57, 16'h9BD1, 16'hB595, 16'hD6DA, 16'hD699, 16'hCE59, 16'hE71C, 16'hFFDF, 16'hFF9E, 16'hEF1C, 16'hDEDB, 16'hDE9A, 16'hDE9A, 16'hD618, 16'hCCD4, 16'hDD14,
        16'hDD55, 16'hDD55, 16'hDD55, 16'hDD55, 16'hDD55, 16'hDD15, 16'hE556, 16'hE556, 16'h7A4A, 16'hE6DC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hA492, 16'h7B0C, 16'h834D, 16'h728A, 16'h934E, 16'hC514, 16'hCD56, 16'hE65A, 16'hE65A,
        16'hDE19, 16'hDE19, 16'hE65A, 16'hDE19, 16'hCD56, 16'hD5D8, 16'hDDD8, 16'hCD56, 16'hBCD4, 16'hB4D3, 16'hB4D3, 16'hBD15, 16'hAC52, 16'hB4D3, 16'hC515, 16'hBD14, 16'hB4D4, 16'hB4D3, 16'hBCD4, 16'hB4D3, 16'hBCD4, 16'hC555, 16'hCD56, 16'hC555, 16'hC556, 16'hC596, 16'hC596, 16'hD618, 16'hD5D7, 16'hC555, 16'hC555, 16'hCD96, 16'hBCD4, 16'hB4D3, 16'hA410, 16'hAC10, 16'h934E, 16'h934D, 16'h934D, 16'h82CB, 16'h8B0C, 16'h8ACB, 16'h934E, 16'hB452, 16'hAC51, 16'hAC51, 16'hC555, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hEE9C, 16'hDE19, 16'hE61A, 16'hEE9B, 16'hEE9B, 16'hBD15, 16'hAC53, 16'hBCD5, 16'hC516, 16'hCD56, 16'hC556, 16'hC556, 16'hCD56, 16'hC516, 16'hC515, 16'hD597, 16'hCD57, 16'hCD97, 16'hC515, 16'hC556, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE1A, 16'hC516, 16'hC515, 16'hBCD5, 16'hCD98, 16'hDE19, 16'hCD97, 16'hCD97, 16'hD5D8, 16'hDE1A, 16'hDE1A, 16'hDE5A, 16'hDE19, 16'hE65A, 16'hDE19, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hDE19, 16'hDE19, 16'hDE5A, 16'hE65A, 16'hE65A, 16'hCD97, 16'hC516,
        16'hC556, 16'hBD15, 16'hCD97, 16'hE65A, 16'hDE19, 16'hDDD9, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hE69B, 16'hE65B, 16'hD598, 16'hB493, 16'hB4D4, 16'hC516, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD57, 16'hC557, 16'hC556, 16'hCD57, 16'hC557, 16'hC556, 16'hC556, 16'hC557, 16'hC556, 16'hC556, 16'hC557, 16'hCD57, 16'h9BD0, 16'hB514, 16'hDEDA, 16'hD699, 16'hD699, 16'hE71C, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF79E, 16'hE6DB, 16'hD69A, 16'hDE9A, 16'hD5D7, 16'hD515, 16'hDD55, 16'hDD55, 16'hDD55, 16'hDD15, 16'hDD15, 16'hDD15, 16'hE556, 16'hD4D4, 16'h6186, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h6249, 16'h000, 16'h4042, 16'h4904, 16'h4883, 16'h6A4A, 16'h938F, 16'hCD56, 16'hE61A, 16'hEE5A, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hF69C, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF71C, 16'hF71D, 16'hEEDC, 16'hEF1C, 16'hEF1C, 16'hEEDC, 16'hEEDC, 16'hF71D, 16'hF71C, 16'hEEDC, 16'hEF1C, 16'hEEDC, 16'hEF1D, 16'hF71D, 16'hF71D, 16'hEF1C, 16'hF71C, 16'hF75D, 16'hEF1C, 16'hF75D, 16'hEF1C, 16'hF75D, 16'hEF1C, 16'hF75D, 16'hF75E, 16'hF79E, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hEEDC, 16'hE61A, 16'hDE19, 16'hE65A, 16'hEE9B, 16'hDE19, 16'hB492, 16'hB493, 16'hC516, 16'hC516, 16'hC515, 16'hC515, 16'hC556, 16'hCD56, 16'hCD56, 16'hBCD5, 16'hD5D8, 16'hD598, 16'hD598, 16'hCD56, 16'hCD57, 16'hE65B, 16'hE69B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hCD56, 16'hC516, 16'hC515, 16'hD5D8, 16'hDE1A, 16'hCD97, 16'hCD97, 16'hD5D8, 16'hDE1A, 16'hDE1A, 16'hE65A, 16'hD5D8, 16'hDE19, 16'hE65B, 16'hDE5A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE1A, 16'hE65A, 16'hE65A, 16'hDE5A, 16'hE65A, 16'hE65A, 16'hD5D8, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hDE1A, 16'hDE19, 16'hCD97, 16'hE69B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE69B, 16'hDE5A, 16'hCD97, 16'hBD15, 16'hC556, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD57, 16'hCD57, 16'hCD57, 16'hC557, 16'hC557, 16'hC556, 16'hCD57, 16'hC557, 16'hC556, 16'hC556, 16'hC557, 16'hC557, 16'hC556, 16'hCD57, 16'h9C11, 16'hAD14, 16'hDE9A, 16'hD699, 16'hD69A,
        16'hEF5D, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF75D, 16'hDEDA, 16'hDE99, 16'hDDD7, 16'hDD55, 16'hDD55, 16'hDD55, 16'hDD15, 16'hE515, 16'hDD15, 16'hE556, 16'hC451, 16'h7B0C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h7B4D, 16'h6186, 16'hABCF, 16'hB3D0, 16'hAB8F, 16'h7A8A, 16'h5186, 16'h51C7, 16'h8B8F, 16'hAC93, 16'hB493, 16'hB493, 16'hB493, 16'hB494, 16'hBC94, 16'hBCD4, 16'hC515, 16'hCD56, 16'hCD57, 16'hCD97, 16'hCD98, 16'hDDD9, 16'hDE19, 16'hDE1A, 16'hDE1A, 16'hE61A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65B, 16'hEE9B, 16'hEE9B, 16'hEEDC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF71D, 16'hE65A, 16'hDE19, 16'hDE1A, 16'hE65A, 16'hE61A, 16'hCD97, 16'hA452, 16'hB494, 16'hC515, 16'hBD15, 16'hC516, 16'hC516, 16'hC516, 16'hC556, 16'hCD97, 16'hBCD4, 16'hCD57, 16'hD5D9, 16'hD5D8, 16'hD598, 16'hCD97, 16'hDE5A, 16'hE69B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65A, 16'hCD97, 16'hC556, 16'hC556, 16'hDE19, 16'hE65A, 16'hD5D8, 16'hCD97, 16'hD598, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hCD98,
        16'hE65B, 16'hE69B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65B, 16'hE65B, 16'hE65B, 16'hD5D9, 16'hCD97, 16'hCD97, 16'hCD57, 16'hC556, 16'hE65A, 16'hDE1A, 16'hCD56, 16'hDE5A, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hDE1A, 16'hCD97, 16'hCD57, 16'hCD98, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD57, 16'hCD57, 16'hCD57, 16'hC556, 16'hCD57, 16'hCD57, 16'hC556, 16'hC557, 16'hC557, 16'hCD57, 16'hCD57, 16'h93D0, 16'hAD14, 16'hD6DA, 16'hCE99, 16'hD69A, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hE6DB, 16'hD618, 16'hDD55, 16'hE555, 16'hDD15, 16'hDD15, 16'hE555, 16'hE556, 16'hE596, 16'hA30D, 16'hA492, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9C51, 16'h69C7, 16'hC452, 16'hC452, 16'hC452, 16'hC451, 16'hAB8F, 16'h828B, 16'h59C7, 16'h730C, 16'hA493, 16'hBD15, 16'hB4D4, 16'hB4D4, 16'hBCD4, 16'hB4D4, 16'hB4D5, 16'hBCD5, 16'hB4D4, 16'hB4D4, 16'hB4D4, 16'hB494, 16'hB494, 16'hB494, 16'hB4D4, 16'hB494, 16'hBC94, 16'hB494, 16'hB494, 16'hBC94, 16'hBCD5, 16'hBC94, 16'hBC94, 16'hBC94, 16'hBC94, 16'hBCD4, 16'hBC94, 16'hB494, 16'hBC94, 16'hBC94, 16'hBC94,
        16'hBC94, 16'hBC94, 16'hC494, 16'hBC94, 16'hC4D4, 16'hCD15, 16'hCD16, 16'hD556, 16'hD597, 16'hDDD8, 16'hE619, 16'hDE19, 16'hE619, 16'hE619, 16'hE65A, 16'hDE1A, 16'hE61A, 16'hE65A, 16'hEE5B, 16'hDE19, 16'hCD57, 16'hC515, 16'hBCD4, 16'hC516, 16'hC515, 16'hC556, 16'hC556, 16'hCD56, 16'hCD57, 16'hD597, 16'hCD56, 16'hBCD4, 16'hDDD9, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hDE5A, 16'hE69B, 16'hE65B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65A, 16'hCD97, 16'hCD56, 16'hCD56, 16'hDE19, 16'hE65A, 16'hDE19, 16'hCD97, 16'hD598, 16'hE65A, 16'hE65B, 16'hE65A, 16'hEE9B, 16'hD5D8, 16'hD5D8, 16'hEE9B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65A, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE69B, 16'hE65B, 16'hEE9B, 16'hDE19, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hE65B, 16'hDE1A, 16'hC516, 16'hDE19, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hDE19, 16'hD5D8, 16'hD5D8, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD57, 16'hCD57, 16'hC556, 16'hCD57,
        16'hCD57, 16'hC557, 16'hC557, 16'hC557, 16'hCD57, 16'h93D0, 16'hAD13, 16'hDED9, 16'hCE99, 16'hD699, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hE69B, 16'hD596, 16'hDD55, 16'hDD15, 16'hDD15, 16'hDD55, 16'hE555, 16'hE556, 16'h8A4A, 16'hB555, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD55, 16'h5800, 16'hBC11, 16'hC452, 16'hC451, 16'hC451, 16'hC452, 16'hC452, 16'hABCF, 16'h7A49, 16'h6187, 16'h93CF, 16'hB4D5, 16'hBCD5, 16'hBCD5, 16'hBCD5, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD16, 16'hBD15, 16'hBD15, 16'hBD16, 16'hBD15, 16'hBD16, 16'hBD16, 16'hBD16, 16'hC516, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC515, 16'hBCD4, 16'hBC93, 16'hC4D4, 16'hBCD4, 16'hC515, 16'hDDD8, 16'hE61A, 16'hE65A, 16'hE65A, 16'hEE5B, 16'hD5D8, 16'hC516, 16'hD5D8, 16'hBCD4, 16'hC515, 16'hCD56, 16'hD597, 16'hD598, 16'hCD97, 16'hCD97, 16'hD598, 16'hD5D8, 16'hBCD4, 16'hCD97, 16'hDE19, 16'hDDD9, 16'hD5D8, 16'hDE1A, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hCD97,
        16'hCD57, 16'hCD57, 16'hDE1A, 16'hE65A, 16'hDE1A, 16'hD597, 16'hD5D8, 16'hE65A, 16'hE69B, 16'hE65B, 16'hE69B, 16'hE65A, 16'hCD56, 16'hE65A, 16'hE69B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hD619, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD98, 16'hEE9B, 16'hE65A, 16'hC515, 16'hDE19, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65A, 16'hE65A, 16'hD5D9, 16'hCD97, 16'hCD97, 16'hCD57, 16'hCD57, 16'hCD97, 16'hCD57, 16'hCD57, 16'hC557, 16'hC557, 16'hCD97, 16'h9C11, 16'hB554, 16'hD699, 16'hD699, 16'hCE58, 16'hEF1C, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hE69A, 16'hD514, 16'hDD15, 16'hDD55, 16'hDD15, 16'hE555, 16'hDD15, 16'h68C4, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h5800, 16'hB3D0, 16'hC452, 16'hC451, 16'hC451, 16'hC452, 16'hC452, 16'hC452, 16'hC451, 16'hA34E, 16'h7187, 16'h728A, 16'hAC93, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD15, 16'hBD16, 16'hBD16, 16'hBD16, 16'hBD15, 16'hBD16, 16'hC516, 16'hC516, 16'hC556, 16'hC556,
        16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hC516, 16'hC556, 16'hC556, 16'hC556, 16'hC516, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC515, 16'hB4D4, 16'hBCD4, 16'hBD15, 16'hBCD4, 16'hC515, 16'hDE19, 16'hE65A, 16'hE65A, 16'hE65A, 16'hEE5B, 16'hD598, 16'hC516, 16'hE61A, 16'hC515, 16'hC515, 16'hD5D8, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD9, 16'hDDD8, 16'hDE19, 16'hCD57, 16'hB493, 16'hDE19, 16'hDE19, 16'hD5D9, 16'hDE19, 16'hE69B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hE69B, 16'hE65B, 16'hEE9B, 16'hE65B, 16'hD5D8, 16'hCD97, 16'hCD97, 16'hE65A, 16'hE65A, 16'hE65A, 16'hD5D8, 16'hD5D8, 16'hE65A, 16'hE69B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hCD97, 16'hD598, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hD5D8, 16'hCD97, 16'hCD97, 16'hCD97, 16'hDE19, 16'hEE9B, 16'hE65A, 16'hC515, 16'hDE19, 16'hEE9C, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B,
        16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hE65A, 16'hDE19, 16'hD598, 16'hCD97, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD97, 16'h93D0, 16'h6249, 16'hB515, 16'hD69A, 16'hCE99, 16'hDEDB, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hF75E, 16'hF75E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hE65A, 16'hD514, 16'hDD55, 16'hDD15, 16'hE555, 16'hCC93, 16'h61C7, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h6A49, 16'hA34D, 16'hC492, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hBC51, 16'hC452, 16'hC492, 16'hBC11, 16'h8A8B, 16'h6186, 16'h93D0, 16'hC515, 16'hBD16, 16'hBD15, 16'hBD15, 16'hBD16, 16'hBD15, 16'hBD16, 16'hC516, 16'hBD16, 16'hC516, 16'hC516, 16'hC556, 16'hC556, 16'hC516, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC557, 16'hC557, 16'hC556, 16'hC556, 16'hC556, 16'hC516, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'hC556, 16'hE61A, 16'hE65B, 16'hE65A, 16'hE65B, 16'hEE5B, 16'hD598, 16'hCD97, 16'hEE9B, 16'hD598, 16'hBD15, 16'hDE19, 16'hDE1A, 16'hDE5A, 16'hDE1A, 16'hDE19, 16'hE65A, 16'hDE19, 16'hDE19, 16'hBC94, 16'hCD97, 16'hE65A,
        16'hDE19, 16'hDE19, 16'hE65B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hE65B, 16'hD5D8, 16'hCD97, 16'hD598, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE19, 16'hD598, 16'hE65A, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hE65A, 16'hC515, 16'hE65B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hCDD8, 16'hCD97, 16'hD598, 16'hD5D8, 16'hE65A, 16'hEE9B, 16'hE65A, 16'hBCD5, 16'hE65A, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hE65B, 16'hE65A, 16'hE65A, 16'hDE1A, 16'hCD98, 16'hCD97, 16'hCD97, 16'hCD57, 16'hCD57, 16'hC556, 16'h93D0, 16'h93D0, 16'h5A08, 16'hBDD6, 16'hD699, 16'hDEDB, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hE71C, 16'hDEDB, 16'hEF1C, 16'hF75D, 16'hF75E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hE618, 16'hD514, 16'hDD15, 16'hE556, 16'hB3CF, 16'h8B8E,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDE, 16'h838E, 16'h8249, 16'hC452, 16'hC452, 16'hC451, 16'hBC51, 16'hC451, 16'hC451, 16'hC452, 16'hC452, 16'hC492, 16'hCC92, 16'hAB8E, 16'h6904, 16'h7B0D, 16'hBD15,
        16'hC516, 16'hBD15, 16'hBD16, 16'hBD15, 16'hBD16, 16'hC516, 16'hC516, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC557, 16'hC556, 16'hC557, 16'hC556, 16'hCD57, 16'hCD57, 16'hC557, 16'hCD57, 16'hCD56, 16'hC556, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hB4D4, 16'hCD57, 16'hE65B, 16'hE69B, 16'hE65A, 16'hEE9B, 16'hE65B, 16'hD5D8, 16'hD5D8, 16'hEE5B, 16'hE61A, 16'hC556, 16'hDE19, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE5A, 16'hE65A, 16'hDE5A, 16'hE65A, 16'hD598, 16'hAC52, 16'hE61A, 16'hDE1A, 16'hDE1A, 16'hE65A, 16'hE69B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hE65B, 16'hDDD9, 16'hD5D8, 16'hD5D8, 16'hE65B, 16'hE69B, 16'hE65B, 16'hE65A, 16'hDDD8, 16'hE61A, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hEE9C, 16'hD597, 16'hD5D9, 16'hEE9C, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hCD97, 16'hD5D8, 16'hCD98,
        16'hDE19, 16'hEE9B, 16'hEE9B, 16'hE61A, 16'hBCD4, 16'hEE9A, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE1A, 16'hCD97, 16'hCD57, 16'hCD57, 16'hCD57, 16'hC516, 16'hC556, 16'hAC52, 16'hC5D7, 16'hE6DB, 16'hE71B, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hEF1C, 16'hD69A, 16'hD69A, 16'hD699, 16'hD6DA, 16'hD6DA, 16'hD6DA, 16'hDE99, 16'hDE17, 16'hD514, 16'hDD14, 16'hE556, 16'h8A8A, 16'hB514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB554, 16'h5000, 16'hBC11, 16'hC452, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hCC52, 16'hCC92, 16'hBC11, 16'h8209, 16'h6A49, 16'hB493, 16'hC556, 16'hBD15, 16'hC516, 16'hC556, 16'hBD16, 16'hC556, 16'hC516, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC557, 16'hC556, 16'hC556, 16'hCD57, 16'hC556, 16'hC556, 16'hC557, 16'hC556, 16'hCD57, 16'hCD57, 16'hCD57, 16'hC557, 16'hCD57, 16'hCD97, 16'hCD56, 16'hBD15, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hD5D8, 16'hE65B, 16'hE65B, 16'hE65A, 16'hE69B, 16'hE65A, 16'hCD97, 16'hDE19, 16'hE65B, 16'hE65A, 16'hD597, 16'hDDD9,
        16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE5A, 16'hE69B, 16'hCD56, 16'hCD57, 16'hE65A, 16'hDE19, 16'hDE5A, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hDE19, 16'hD5D8, 16'hDDD8, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE65B, 16'hDE19, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hEE9C, 16'hE65A, 16'hCD57, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hDE19, 16'hCD98, 16'hD5D8, 16'hD5D9, 16'hE65B, 16'hE69B, 16'hEE9C, 16'hD5D9, 16'hC515, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE65B, 16'hDE19, 16'hC556, 16'hCD97, 16'hCD97, 16'hCD97, 16'h938F, 16'h7B0C, 16'hCDD8, 16'hD699, 16'hF75D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hF75D,
        16'hDE9A, 16'hD659, 16'hD618, 16'hCDD7, 16'hCD96, 16'hD595, 16'hD514, 16'hD514, 16'hDD15, 16'hD4D4, 16'h6946, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDA, 16'h4000, 16'hABCF, 16'hCC92,
        16'hC451, 16'hC452, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC452, 16'hCC92, 16'hC452, 16'h92CB, 16'h50C3, 16'hA452, 16'hC557, 16'hC516, 16'hBD16, 16'hC516, 16'hC516, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC557, 16'hC556, 16'hCD57, 16'hCD57, 16'hCD57, 16'hC557, 16'hCD57, 16'hCD57, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hC556, 16'hBCD4, 16'hBCD4, 16'hBCD4, 16'hD5D8, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hCD97, 16'hDE19, 16'hE65B, 16'hE65A, 16'hDE19, 16'hD598, 16'hE65A, 16'hE65B, 16'hE65A, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65B, 16'hE61A, 16'hB452, 16'hDE19, 16'hDE5A, 16'hDE5A, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hE65B, 16'hDE19, 16'hD5D8, 16'hDE19, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hD597, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B,
        16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hD5D9, 16'hD5D8, 16'hD619, 16'hE65A, 16'hEE9B, 16'hE65B, 16'hEE9C, 16'hCD57, 16'hCD57, 16'hEE9C, 16'hE69B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hE69B, 16'hE65B, 16'hE69B, 16'hE65B, 16'hE65A, 16'hE65B, 16'hE69B, 16'hD5D8, 16'hBD15, 16'hCD97, 16'h93D0, 16'h5187, 16'hAC93, 16'hA493, 16'hCE58, 16'hE71C, 16'hEF1C, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hF79E, 16'hD618, 16'hCC92, 16'hCC52, 16'hCC92, 16'hD4D3, 16'hD4D4, 16'hD514, 16'hDD15, 16'hBC11, 16'h7B0C, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h8B8E, 16'h8ACB, 16'hD514, 16'hC492, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC452, 16'hCC92, 16'hCC92, 16'hAB8E, 16'h6987, 16'h9BD0, 16'hC516, 16'hC556, 16'hC516, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC557, 16'hC557, 16'hC556, 16'hC557, 16'hC557, 16'hC556, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD97, 16'hCD57, 16'hCD57, 16'hCD97, 16'hCD97, 16'hCD97, 16'hC515, 16'hBD15, 16'hBD15, 16'hD5D8, 16'hE69B,
        16'hE69B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hCD57, 16'hD619, 16'hE69B, 16'hE65A, 16'hE65A, 16'hD5D8, 16'hDE1A, 16'hEE5B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65B, 16'hE65B, 16'hEE9C, 16'hCD16, 16'hB493, 16'hEE9B, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hDE19, 16'hDE19, 16'hDE19, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hDE1A, 16'hDE19, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hD5D9, 16'hD619, 16'hE65A, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hC515, 16'hDDD8, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE69B, 16'hCD97, 16'hC516, 16'hBCD4, 16'h6A4A, 16'hBD55, 16'hEF1C, 16'hE6DB, 16'hE6DB, 16'hE6DB,
        16'hE71C, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF5E, 16'hD556, 16'hCC52, 16'hD4D3, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hDD15, 16'h92CB, 16'hA493, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD14, 16'h5882, 16'hD514, 16'hD514, 16'hCCD3, 16'hC492, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC452, 16'hC452, 16'hC452, 16'hC452, 16'hB3D0, 16'h7187, 16'h82CC, 16'hBD15, 16'hC556, 16'hC516, 16'hC516, 16'hC556, 16'hC556, 16'hC556, 16'hC557, 16'hC557, 16'hC556, 16'hC557, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD97, 16'hCD57, 16'hCD97, 16'hCD97, 16'hCD97, 16'hC556, 16'hC515, 16'hD598, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hC556, 16'hD597, 16'hE69B, 16'hE65B, 16'hE65B, 16'hDE19, 16'hD5D8, 16'hEE5B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hAB90, 16'hDE19, 16'hE69B, 16'hDE5A, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hDE1A, 16'hDE19, 16'hDE1A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE65A,
        16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hDDD9, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hDE19, 16'hE65A, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hC515, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE69B, 16'hEE9B, 16'hBD15, 16'h8B4D, 16'h728B, 16'h9C51, 16'hE6DC, 16'hE6DB, 16'hE6DB, 16'hE71C, 16'hE6DB, 16'hE6DC, 16'hF75D, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hF75D, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hCD14, 16'hCC93, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'h6945, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h4841, 16'hC452, 16'hE556, 16'hDD55, 16'hDD15, 16'hCCD3, 16'hC451, 16'hC451, 16'hC451, 16'hC451, 16'hC452, 16'hC452, 16'hC452, 16'hC452, 16'hC451, 16'hC492, 16'hBD14, 16'h9C10, 16'h724A, 16'hAC53, 16'hCD57, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC557, 16'hC557, 16'hC557, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD57,
        16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD98, 16'hCD97, 16'hC556, 16'hD598, 16'hE65B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hCD57, 16'hC556, 16'hE69B, 16'hE65B, 16'hE69B, 16'hE65A, 16'hD5D8, 16'hE61A, 16'hEE9B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hEE9C, 16'hDD98, 16'hB451, 16'hF71D, 16'hE65A, 16'hE65A, 16'hE69B, 16'hEE9C, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE65A, 16'hDE1A, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hE61A, 16'hE65A, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hEE9C, 16'hD5D8, 16'hCD56, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B,
        16'hE69B, 16'hE69B, 16'hE65B, 16'hE69B, 16'hE65A, 16'h7B0D, 16'h834E, 16'hDE19, 16'hDEDB, 16'hE6DB, 16'hE6DB, 16'hE6DB, 16'hE6DB, 16'hE6DC, 16'hE6DB, 16'hEF1C, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hF75E, 16'hDE9B, 16'hE6DB, 16'hEF1C, 16'hFF5E, 16'hFF9F, 16'hFFDF, 16'hEEDB, 16'hCC93, 16'hD4D3, 16'hD4D4, 16'hDD14, 16'hABCF, 16'h7B0B, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h838E, 16'h92CC, 16'hE556, 16'hDD56, 16'hDD55, 16'hDD15, 16'hD514, 16'hCC92, 16'hC452, 16'hC452, 16'hC451, 16'hC451, 16'hCC92, 16'hCC51, 16'hC492, 16'hC556, 16'hC5D7, 16'hC5D7, 16'hAD13, 16'h7B0C, 16'hA411, 16'hC556, 16'hCD57, 16'hC556, 16'hC556, 16'hC557, 16'hC557, 16'hC557, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD97, 16'hCD97, 16'hCD57, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hD5D8, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hEEDC, 16'hD597, 16'hBCD4, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hDE19, 16'hDE19, 16'hEE9B, 16'hE65B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hF6DC, 16'hB3D1, 16'hD5D7, 16'hFF5E, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B,
        16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE65A, 16'hE65A, 16'hE65B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hE65B, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hDE19, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hC515, 16'hD5D8, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hEE9B, 16'hEE9B, 16'h7B0C, 16'hB4D4, 16'hEF1C, 16'hE71C, 16'hEF1D, 16'hEF1C, 16'hE6DB, 16'hE6DB, 16'hE6DB, 16'hE6DB, 16'hE6DB, 16'hEF5D, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hD659, 16'hCD96, 16'hB451, 16'hD596, 16'hE659, 16'hEE9A, 16'hD515, 16'hCC92, 16'hD4D3, 16'hDD14, 16'h7186, 16'hC596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD658, 16'h5800, 16'hD514, 16'hE596, 16'hDD55, 16'hDD55, 16'hDD56, 16'hDD55, 16'hCCD3, 16'hC452, 16'hC451, 16'hC451, 16'hC452, 16'hC4D3, 16'hBD95, 16'hC5D7, 16'hCE19, 16'hD69A, 16'hD699, 16'hC5D7, 16'h9C10, 16'h938F,
        16'hB494, 16'hC557, 16'hC557, 16'hC557, 16'hC556, 16'hC557, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hD5D8, 16'hE65B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hDE19, 16'hB453, 16'hE65A, 16'hE69B, 16'hE65B, 16'hE65B, 16'hE65A, 16'hDE19, 16'hE65B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hE61A, 16'h9ACC, 16'hF75D, 16'hF71D, 16'hE61A, 16'hE65A, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hE65A, 16'hE69B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hDE19, 16'hE65B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hEEDC,
        16'hDE19, 16'hC4D5, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hE69B, 16'hE65B, 16'hE69B, 16'hE65B, 16'hE65B, 16'hEE9B, 16'hD5D8, 16'h4904, 16'hCDD7, 16'hE6DB, 16'hF75D, 16'hFFDF, 16'hFF9E, 16'hF75D, 16'hEF1C, 16'hEF1C, 16'hE6DC, 16'hE6DB, 16'hE6DC, 16'hF75D, 16'hFF9E, 16'hFF9F, 16'hEF1C, 16'hDE59, 16'hBC51, 16'hBBCF, 16'hC411, 16'hC451, 16'hCC92, 16'hCC92, 16'hD4D4, 16'hB3CF, 16'h5987, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h72CB, 16'hB3D0, 16'hE597, 16'hDD56, 16'hDD56, 16'hDD56, 16'hDD56, 16'hDD55, 16'hD4D4, 16'hCC92, 16'hCC51, 16'hC492, 16'hC596, 16'hCE18, 16'hDE9B, 16'hE6DC, 16'hE71C, 16'hE6DB, 16'hDEDB, 16'hCE18, 16'hACD3, 16'h7B0C, 16'h9C11, 16'hBD56, 16'hCD97, 16'hC557, 16'hCD97, 16'hCD57, 16'hCD57, 16'hC557, 16'hCD57, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hD598, 16'hE65A, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65A, 16'hB453, 16'hDE19, 16'hEE9B, 16'hE69B, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hD556, 16'hA3D0, 16'hFFDF,
        16'hEEDC, 16'hE61A, 16'hE65B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hE61A, 16'hDDD9, 16'hEEDC, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hC4D5, 16'hD597, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hEE9B, 16'hB493, 16'h7B0D, 16'hE69A, 16'hDE9A, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hF75E, 16'hF75D, 16'hEF1D, 16'hEF1D, 16'hF75E, 16'hFF9E, 16'hEF1D, 16'hDE59, 16'hC453, 16'hC412, 16'hCC93, 16'hCC92, 16'hCC93, 16'hD4D3, 16'h60C4,
        16'hBD15, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB555, 16'h79C8, 16'hE556, 16'hDD96, 16'hDD56, 16'hDD56, 16'hDD56, 16'hDD56, 16'hDD55,
        16'hD4D4, 16'hD513, 16'hDE18, 16'hE71B, 16'hEF1D, 16'hF75D, 16'hEF1C, 16'hE6DB, 16'hE6DB, 16'hE71C, 16'hDE9A, 16'hCE18, 16'hC596, 16'hA451, 16'h7B0C, 16'hA453, 16'hCD57, 16'hCD57, 16'hCD97, 16'hCD57, 16'hCD57, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hD598, 16'hCD97, 16'hDE19, 16'hE69B, 16'hE65B, 16'hE69B, 16'hE69B, 16'hEE9C, 16'hBCD5, 16'hD597, 16'hEE9B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE69B, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hA34E, 16'hCD96, 16'hFFDF, 16'hEEDC, 16'hE61A, 16'hE65B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE5B, 16'hCD57, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B,
        16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hDE19, 16'hBC93, 16'hDE1A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hEE5B, 16'h7ACC, 16'hBD55, 16'hDE9B, 16'hD659, 16'hDE9B, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hF75E, 16'hEEDB, 16'hD556, 16'hC492, 16'hC451, 16'hC451, 16'h9B0C, 16'h3000, 16'h938E, 16'h8BCF, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h5945, 16'hC492, 16'hE597, 16'hDD56, 16'hE556, 16'hE556, 16'hDD56, 16'hDD56, 16'hD514, 16'hDD97, 16'hEEDB, 16'hEEDC, 16'hEEDC, 16'hEEDB, 16'hE69B, 16'hDEDB, 16'hE6DB, 16'hE6DB, 16'hEF1C, 16'hF75D, 16'hEF1C, 16'hCE18, 16'hB514, 16'h8B8E, 16'h9BD0, 16'hC556, 16'hCD97, 16'hCD97, 16'hCD57, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hD598, 16'hD5D9, 16'hE65A, 16'hE65B, 16'hE65B, 16'hE65B, 16'hEE9B, 16'hD597, 16'hC4D4, 16'hF6DC, 16'hE65A, 16'hEE9B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hEE9B,
        16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEEDC, 16'hE65A, 16'h924A, 16'hEF1C, 16'hFFDF, 16'hEE9C, 16'hE65A, 16'hE69B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hD556, 16'hE619, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hC4D4, 16'hCD56, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hEE9B, 16'hC556, 16'h728A, 16'hDE59, 16'hDE9A, 16'hD659, 16'hD659, 16'hDE9A, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E,
        16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hF75D, 16'hEEDC, 16'hE65A, 16'hD596, 16'hBCD3, 16'hBCD3, 16'h4000, 16'h9411, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA451, 16'h928C, 16'hE597, 16'hDD96, 16'hE596, 16'hDD56, 16'hE556, 16'hE556, 16'hDD14, 16'hD4D3, 16'hCC93, 16'hCC93, 16'hCC52, 16'hBC10, 16'hD5D7, 16'hDE9A, 16'hE71C, 16'hF75D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hEF1D, 16'hD69A, 16'hD618, 16'h938F, 16'h830D, 16'hB4D4, 16'hC556, 16'hCD57, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hD5D8, 16'hD5D8, 16'hE65A, 16'hE69B, 16'hE65A, 16'hE65B, 16'hE69B, 16'hEE5B, 16'hABD1, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hE69B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEEDC, 16'hCCD5, 16'h92CC, 16'hFF9F, 16'hFFDF, 16'hEE9C, 16'hE61A, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B,
        16'hF6DC, 16'hDDD8, 16'hCD56, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hDDD9, 16'hB453, 16'hDE19, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hE65B, 16'hEE9B, 16'h9BCF, 16'h9410, 16'hDE9A, 16'hDE9A, 16'hEF1C, 16'hF75D, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hF79E, 16'hF75E, 16'hF75E, 16'hF79E, 16'hF75E, 16'hFF5D, 16'hC596, 16'h830C, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h6000, 16'hD514, 16'hE597, 16'hE556, 16'hE556, 16'hE556, 16'hE556, 16'hE556, 16'hDD15, 16'hDD15, 16'hDCD4, 16'hC38F, 16'hC452, 16'hE659, 16'hF71D, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hEF1D, 16'hC596, 16'h728A, 16'h82CC, 16'hB4D4, 16'hC556, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hC556, 16'hD5D8, 16'hE65A, 16'hE65A, 16'hEEDC, 16'hE65A, 16'hE65B, 16'hE65A,
        16'hEE9C, 16'hCCD5, 16'hD597, 16'hFF1D, 16'hE65A, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF69B, 16'hAB4E, 16'hC493, 16'hFFDF, 16'hFFDF, 16'hEE9C, 16'hE61A, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hEE5A, 16'hC493, 16'hEE5A, 16'hEEDC, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hBC94, 16'hC516, 16'hE65B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hE69B, 16'hE69B, 16'hE65B,
        16'hE69B, 16'hE619, 16'h61C7, 16'hC596, 16'hE6DB, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hF79E, 16'hF75E, 16'hFF9E, 16'hF79E, 16'hF75D, 16'hCDD8, 16'h4000, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h93CF, 16'h9ACC, 16'hED57, 16'hE556, 16'hE556, 16'hE556, 16'hE556, 16'hE556, 16'hE557, 16'hE597, 16'hDD15, 16'hCCD3, 16'hEE9A, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hEF1D, 16'hD659, 16'hCE18, 16'hACD3, 16'hA452, 16'hAC92, 16'hAC93, 16'hC556, 16'hCD97, 16'hCD97, 16'hCD57, 16'hD5D8, 16'hF69C, 16'hF6DC, 16'hFF9F, 16'hEE9C, 16'hE65A, 16'hE65B, 16'hE69B, 16'hE65A, 16'hA38F, 16'hF75D, 16'hEEDC, 16'hE65B, 16'hE65B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEEDC, 16'hE61A, 16'h9107, 16'hE5D9, 16'hFFDF, 16'hFFDF, 16'hEE9C, 16'hE61A, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C,
        16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hC494, 16'hDD97, 16'hF6DC, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hDD98, 16'hB452, 16'hDDD9, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hEE9C, 16'hB493, 16'h834D, 16'hDE9A, 16'hE71C, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hF75E, 16'hF75D, 16'hEF1C, 16'hDE9A, 16'hACD3, 16'h4000, 16'hBD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h5800, 16'hCC93, 16'hE557, 16'hE556, 16'hE556, 16'hE556, 16'hE556, 16'hE556, 16'hE556, 16'hDD15, 16'hEE9A, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hDE9B, 16'hDE9A, 16'hDE9A, 16'hE6DB, 16'hDE19, 16'h9BD0, 16'hA452,
        16'hCD97, 16'hB493, 16'hC4D5, 16'hDDD9, 16'hF6DD, 16'hFF5E, 16'hFFDF, 16'hFF9F, 16'hEE5B, 16'hEE9B, 16'hE65A, 16'hEE9B, 16'hBC93, 16'hC515, 16'hFF9E, 16'hE65B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hDD57, 16'hA20A, 16'hF69B, 16'hFFDF, 16'hFF9F, 16'hEE9C, 16'hE65A, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hCD16, 16'hC494, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hE65A, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE5B, 16'hBC94, 16'hCD15, 16'hE65A, 16'hEE9B,
        16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hE65B, 16'hE69B, 16'hEE5A, 16'h724A, 16'hB515, 16'hDEDB, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hF75E, 16'hFF9F, 16'hFF9E, 16'hF79E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hF75D, 16'hD619, 16'h72CB, 16'h000, 16'h7B4D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h8B8E, 16'h930C, 16'hE596, 16'hE556, 16'hE556, 16'hE556, 16'hE556, 16'hE556, 16'hDD15, 16'hEE5A, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9F, 16'hE69B, 16'h9C10, 16'hAC92, 16'hD5D8, 16'hAC12, 16'hB412, 16'hF65B, 16'hFF1E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF5F, 16'hFF1E, 16'hEEDC, 16'hEE9B, 16'hE619, 16'h9ACD, 16'hF71D, 16'hF71D, 16'hE65A, 16'hE65B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hE65B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hBC52, 16'hBB0F, 16'hF71D, 16'hFFDF, 16'hFF9F, 16'hEE9C, 16'hEE5A, 16'hF6DC, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEE9C,
        16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hF69C, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEE9C, 16'hEEDC, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hE5D9, 16'hB3D1, 16'hE65A, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF69C, 16'hE61A, 16'hEE5B, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hD597, 16'hB453, 16'hE619, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hEE9B, 16'hBCD4, 16'h830C, 16'hDE9A, 16'hE6DB, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hE71C, 16'hF75D, 16'hFF9E, 16'hEF1C, 16'hE6DB, 16'hEF1C, 16'hEF1C, 16'hEF1C, 16'hEF1C, 16'hD618, 16'hAC51, 16'h72CB, 16'h93CF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h5000, 16'hCCD4, 16'hE557, 16'hE556, 16'hE556, 16'hE556, 16'hDD56, 16'hE618, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hCE18, 16'hC597, 16'hDE59, 16'hAC52, 16'hA34F, 16'hFEDD, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hF71D, 16'hEEDC, 16'hB452, 16'hBCD4, 16'hFFDF, 16'hEE9B, 16'hE65B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hE65B, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE5B, 16'hAB4F, 16'hCC12, 16'hFF5E, 16'hFFDF, 16'hFF9F, 16'hEE5B, 16'hEE5A, 16'hF6DC, 16'hEE9C, 16'hF6DC, 16'hF6DC, 16'hF69C, 16'hF69C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hEE9C, 16'hF69C, 16'hF69C, 16'hF69C, 16'hF69C, 16'hF69C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hE65B, 16'hEE9C, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEE9B, 16'hB3D1, 16'hDD98, 16'hF6DC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hE65A, 16'hE619, 16'hEEDC, 16'hEE9B, 16'hEE9C, 16'hEE9C,
        16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE61A, 16'hB452, 16'hD557, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hE69B, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hE69B, 16'hE65B, 16'hE65B, 16'hE69B, 16'hE65A, 16'h82CC, 16'hC556, 16'hDE9A, 16'hEF1C, 16'hFF9F, 16'hFF9F, 16'hE71C, 16'hDE9A, 16'hEF1C, 16'hEF1C, 16'hD659, 16'hDE5A, 16'hDE5A, 16'hDE9A, 16'hDE5A, 16'hD659, 16'hC555, 16'h4103, 16'h838E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA491, 16'h8A4A, 16'hE556, 16'hE556, 16'hE556, 16'hE556, 16'hDD55, 16'hE5D8, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hE659, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hDEDB, 16'hDE9A, 16'hDE9A, 16'hBCD4, 16'h824A, 16'hF6DC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hEE5B, 16'h89C8, 16'hEEDC, 16'hFF9F, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hE5D9, 16'hAACD,
        16'hDD15, 16'hFF9E, 16'hFFDF, 16'hFF5F, 16'hEE5B, 16'hEE5A, 16'hFEDD, 16'hEE9C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF69C, 16'hF69C, 16'hEE9C, 16'hEE9C, 16'hF69C, 16'hF6DC, 16'hEE9B, 16'hE61A, 16'hEE9B, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEE9C, 16'hF6DC, 16'hBC52, 16'hCCD5, 16'hF69C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hEE5B, 16'hD598, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hF75D, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hC4D5, 16'hBC93, 16'hE61A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE65B, 16'hE69B, 16'hE65B, 16'hEE9C, 16'hBCD5, 16'h8B8E, 16'hDE9A, 16'hD65A, 16'hEF1D, 16'hFFDF, 16'hEF1C, 16'hD65A, 16'hDE9A, 16'hDE9B, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hDE5A, 16'hD619, 16'hACD4,
        16'h6A8B, 16'h7B0D, 16'h3882, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D,
        16'h7249, 16'hC452, 16'hE556, 16'hE556, 16'hDD56, 16'hE555, 16'hDD15, 16'hDCD4, 16'hD494, 16'hCC52, 16'hE619, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hE6DB, 16'hE6DB, 16'hE71B, 16'hD618, 16'h7106, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD16, 16'hAC11, 16'hFFDF, 16'hFF9F, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hEE9B, 16'hEE9B, 16'hDE19, 16'hE65B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hF6DC, 16'hCCD4, 16'hC411, 16'hE597, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hF65B, 16'hEE5B, 16'hFEDD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hF69C, 16'hF69C, 16'hF69C, 16'hF6DC, 16'hEE9C, 16'hDE19, 16'hEE5A, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hEEDC, 16'hEE9C, 16'hF69C, 16'hEE9C, 16'hF6DC, 16'hCD15, 16'hB3D1, 16'hF65B, 16'hEEDC, 16'hEEDC,
        16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEEDC, 16'hD598, 16'hDE19, 16'hEE9B, 16'hF71D, 16'hF71D, 16'hEEDC, 16'hFFDF, 16'hF79E, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hDDD8, 16'hABD0, 16'hDD98, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE69B, 16'hE65A, 16'h7ACB, 16'hC597, 16'hDE9B, 16'hDE5A, 16'hEF1D, 16'hEF1C, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hBD96, 16'h5187, 16'hA492, 16'hB515, 16'h4945, 16'h9C51, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD55, 16'h79C7, 16'hE556, 16'hDD56, 16'hDD55, 16'hDD15, 16'hDD15, 16'hDD15, 16'hD493, 16'hE619, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF75D, 16'hF75D, 16'hF75D, 16'hF71D, 16'h9B4E, 16'hCD56, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'h9A8C, 16'hE69A, 16'hFFDF, 16'hFF9F, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hEE9B, 16'hE65A,
        16'hDDD9, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF69C, 16'hBC12, 16'hDD16, 16'hE5D8, 16'hFFDF, 16'hFF9F, 16'hFF1E, 16'hF65B, 16'hF65B, 16'hFEDD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF69C, 16'hEE9C, 16'hF69C, 16'hF69C, 16'hF69C, 16'hF6DC, 16'hF69C, 16'hDDD8, 16'hE61A, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hF6DC, 16'hEE9C, 16'hF6DC, 16'hE5D9, 16'hA30E, 16'hE619, 16'hF6DC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF69C, 16'hEE9C, 16'hF71D, 16'hF6DC, 16'hDDD9, 16'hD597, 16'hEE9B, 16'hF71C, 16'hFFDF, 16'hEE9C, 16'hFF9E, 16'hFFDF, 16'hEEDC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hE65A, 16'hB411, 16'hCD16, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hE65B, 16'hE65B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE65B, 16'hEE9B, 16'hE65B, 16'hE65A, 16'hE69B, 16'hE65B, 16'hEE9B, 16'hAC92, 16'h9C11, 16'hDE9A,
        16'hD65A, 16'hD65A, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hDE5A, 16'hDE5A, 16'hDE9A, 16'hDE9A, 16'hDE5A, 16'hDE5A, 16'h9451, 16'h6249, 16'hACD4, 16'h9C51, 16'h2000, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'h830C, 16'hBC10, 16'hE556, 16'hDD15, 16'hDD15, 16'hE515, 16'hD4D4, 16'hDD97, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hCD56, 16'hAB8F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE19, 16'hAB8F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE619, 16'hE619, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hF69C, 16'hE5D9, 16'hB390, 16'hEDD9, 16'hE5D8, 16'hFFDF, 16'hFF9F, 16'hFF1E, 16'hF65B, 16'hF65B, 16'hFF1D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF69C, 16'hF69C, 16'hEE9C, 16'hF69C, 16'hF69C, 16'hF71D, 16'hF71D, 16'hF69C, 16'hDDD9, 16'hD597, 16'hF69C,
        16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hEE5A, 16'h9ACC, 16'hD557, 16'hF6DC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hFF9F, 16'hF6DD, 16'hEE5B, 16'hCD56, 16'hE65A, 16'hEEDC, 16'hEEDC, 16'hEE9B, 16'hEEDC, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hC4D4, 16'hA3D1, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hEE9B, 16'hEEDC, 16'hE65B, 16'hE65B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hE65B, 16'hE61A, 16'hE65A, 16'hE65B, 16'hE69B, 16'hD5D8, 16'h830D, 16'hCDD8, 16'hD65A, 16'hD65A, 16'hD65A, 16'hD65A, 16'hD659, 16'hD619, 16'hD619, 16'hD619, 16'hD659, 16'hDE5A, 16'hE69B, 16'hD619, 16'h834D, 16'h838F, 16'hBD55, 16'h5186, 16'h9C92, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCDD7, 16'h5000, 16'hD4D4, 16'hDD15, 16'hDD15, 16'hDD15, 16'hDD56, 16'hFF5E, 16'hFFDF, 16'hFF9F, 16'hF75E, 16'hF75D, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF6DC, 16'h9ACB, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5F, 16'hFF5F, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFF9F, 16'hB390, 16'hDDD8, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hDDD9, 16'hE65A, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hF69C, 16'hEE9C, 16'hF69C, 16'hEE9B, 16'hF6DC, 16'hD515, 16'hB412, 16'hEE1A, 16'hE61A, 16'hFFDF, 16'hFF1E, 16'hFF1E, 16'hF65B, 16'hF61A, 16'hFF1D, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hFF1D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9B, 16'hF6DC, 16'hFEDD, 16'hFF5F, 16'hFF5E, 16'hF69C, 16'hE619, 16'hD516, 16'hF69B, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hEEDC, 16'hF69C, 16'hAB8F, 16'hBC94, 16'hF6DC, 16'hEE9C, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DD, 16'hEE9C, 16'hF69C, 16'hD556, 16'hD5D8, 16'hEEDC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hD598, 16'h92CD, 16'hD5D7, 16'hEEDC, 16'hE65B, 16'hF6DC, 16'hF75D, 16'hE69B, 16'hFFDF, 16'hF71D,
        16'hE65B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hEE5B, 16'hE65A, 16'hDE1A, 16'hE65B, 16'hE65B, 16'hEE5B, 16'h938F, 16'hAC92, 16'hD659, 16'hD659, 16'hD659, 16'hDE5A, 16'hD659, 16'hCE19, 16'hCE19, 16'hC597, 16'hA492, 16'hB514, 16'hB514, 16'hBD55, 16'hB514, 16'h6249, 16'hACD3, 16'h9410, 16'h3040, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA492, 16'h8209, 16'hE515, 16'hDD15, 16'hDCD4, 16'hEE19, 16'hEE9B, 16'hE619, 16'hE659, 16'hEEDB, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB411, 16'hCD95, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF6DC, 16'hAB0D, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hD5D8, 16'hEE5B, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hF69C, 16'hBBD1, 16'hCD56, 16'hF5DA, 16'hE65A, 16'hFFDF, 16'hFF1E, 16'hFF1E, 16'hF61B, 16'hEE1A, 16'hFF1D, 16'hF6DC, 16'hF6DD, 16'hFEDD, 16'hFEDD, 16'hFF1D, 16'hF6DC, 16'hF6DC, 16'hFF1D, 16'hF6DC, 16'hF6DC, 16'hFF1D, 16'hFF1D, 16'hFF5E,
        16'hF6DC, 16'hF6DC, 16'hF69C, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hFF1E, 16'hFF1E, 16'hF69C, 16'hE61A, 16'hCCD5, 16'hEE5A, 16'hF6DC, 16'hEEDC, 16'hF69C, 16'hF69C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hBC53, 16'hABD0, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hF69C, 16'hDD98, 16'hCD57, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hA38F, 16'hBC94, 16'hEE9B, 16'hE65B, 16'hEEDC, 16'hFFDF, 16'hEEDB, 16'hF75D, 16'hFF9F, 16'hE69B, 16'hE65B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65A, 16'hDE19, 16'hE65B, 16'hE65A, 16'hE69B, 16'hBD15, 16'h8B4D, 16'hCDD7, 16'hD619, 16'hD659, 16'hD659, 16'hD659, 16'hCE19, 16'hCE18, 16'hCE18, 16'h9C51, 16'h000, 16'h4985, 16'h628A, 16'h6A8A, 16'h6249, 16'h9410, 16'hB4D4, 16'h1800, 16'hB514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h830C, 16'hA34E, 16'hD4D3, 16'hCC52, 16'hCC52, 16'hCCD3, 16'hDDD8, 16'hF71D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE19, 16'h9B4D,
        16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDD57, 16'hC493, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'hEE5B, 16'hEE9B, 16'hE61A, 16'hDDD8, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hF69C, 16'hEE9C, 16'hF65B, 16'hAACE, 16'hE61A, 16'hEDD9, 16'hEE5A, 16'hFF9F, 16'hF6DD, 16'hFF1E, 16'hF65B, 16'hEE5B, 16'hFF1E, 16'hF6DC, 16'hF6DD, 16'hFEDD, 16'hFF1D, 16'hFF5E, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE5B, 16'hEE9B, 16'hF69C, 16'hF69C, 16'hF69C, 16'hF69C, 16'hEE5B, 16'hCCD5, 16'hDDD9, 16'hF6DC, 16'hEE9C, 16'hF69C, 16'hF69C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DD, 16'hD556, 16'h92CC, 16'hE65A, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hE61A, 16'hC515, 16'hE65B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B,
        16'hEE9B, 16'hE69B, 16'hEE9B, 16'hBC93, 16'h9B8F, 16'hE65B, 16'hE69B, 16'hE69B, 16'hEEDC, 16'hEE9B, 16'hE69B, 16'hEE9C, 16'hE69B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE69B, 16'hE65B, 16'hDE19, 16'hDE1A, 16'hE65B, 16'hE65A, 16'hDDD8, 16'h82CC, 16'hBD55, 16'hCE19, 16'hCE19, 16'hCE19, 16'hCE19, 16'hD619, 16'hCE19, 16'hCE18, 16'hCE18, 16'hACD3, 16'h6249, 16'hA492, 16'hB514, 16'hACD3, 16'hACD4, 16'hB515, 16'h628A, 16'h4103, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD14, 16'h5883, 16'hC4D3, 16'hE618, 16'hF6DB, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hA30D, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hBBD1, 16'hE659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hF71D, 16'hF6DC, 16'hDD98, 16'hDDD8, 16'hF71D, 16'hF6DD, 16'hF71D, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hF69C, 16'hF69C, 16'hE5D9, 16'h9A4B, 16'hF6DC, 16'hEDD9, 16'hEE5B, 16'hFF5E, 16'hF69C, 16'hFF1E, 16'hF61B, 16'hEE5B, 16'hFF1E, 16'hF6DC,
        16'hF6DD, 16'hF6DD, 16'hFEDD, 16'hF71D, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE1A, 16'hEE9B, 16'hF6DC, 16'hEE9C, 16'hF69C, 16'hF69C, 16'hF69B, 16'hCD15, 16'hD597, 16'hF6DC, 16'hEE9C, 16'hF69C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hE5D8, 16'h8209, 16'hDDD8, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hC4D5, 16'hDE19, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hEE9C, 16'hCD57, 16'h8ACC, 16'hDE19, 16'hEE9B, 16'hE69B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE69B, 16'hDE1A, 16'hD5D9, 16'hE65A, 16'hDE5A, 16'hE65A, 16'h9BD0, 16'h9410, 16'hD659, 16'hCE18, 16'hCE18, 16'hCE18, 16'hCE18, 16'hCE19, 16'hCE19, 16'hCE18, 16'hD659, 16'hAD14, 16'h59C7, 16'hA493, 16'hB555, 16'hB515, 16'hBD55, 16'h9410, 16'h800, 16'h9410, 16'hFF9E,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h4800, 16'hAC11, 16'hF71C, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD55, 16'hBCD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF69C, 16'hB30D, 16'hFF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hFFDF, 16'hF6DC, 16'hCD15, 16'hE65A, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hEE9B, 16'hEE9C, 16'hF69C, 16'hEE9C, 16'hF6DC, 16'hD556, 16'hAB90, 16'hFF1E, 16'hEDD9, 16'hEE1A, 16'hFF1D, 16'hF69C, 16'hFEDD, 16'hEDDA, 16'hE619, 16'hFEDD, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hE61A, 16'hEE5B, 16'hF69C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF69C, 16'hD557, 16'hCD15, 16'hF69C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hE61A, 16'h8209, 16'hCD56, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B,
        16'hEE9B, 16'hC515, 16'hCD97, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hDDD9, 16'h8ACC, 16'hC556, 16'hEE9B, 16'hE69B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65A, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE65B, 16'hE65A, 16'hD5D8, 16'hDE5A, 16'hE65A, 16'hE65A, 16'hC516, 16'h728A, 16'hC5D6, 16'hCE19, 16'hCE18, 16'hCE18, 16'hCE18, 16'hCE18, 16'hCDD8, 16'hC5D7, 16'hCDD8, 16'hDE5A, 16'hACD3, 16'h6289, 16'hA492, 16'hB514, 16'hBD55, 16'hBD55, 16'h5A49, 16'h6A4A, 16'hC596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hA410, 16'h8B0C, 16'hC555, 16'hEE9B, 16'hF75D, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hE69A, 16'h8A49, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF1E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hE557, 16'hCC53, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF6DC, 16'hFF9E, 16'hE61A, 16'hCD16, 16'hEE5B, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEE9B, 16'hEE9C, 16'hF69C, 16'hEE9C, 16'hF6DC,
        16'hBC52, 16'hBC93, 16'hFF5E, 16'hE598, 16'hE619, 16'hF6DC, 16'hF69C, 16'hFEDD, 16'hE5D9, 16'hE5D8, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF69C, 16'hE61A, 16'hE65A, 16'hF69C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hF69C, 16'hDD98, 16'hC493, 16'hEE5B, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5A, 16'h828A, 16'hB493, 16'hE65A, 16'hE65B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE9C, 16'hD597, 16'hC4D5, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hE61A, 16'h9B4F, 16'hAC52, 16'hEE9B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65B, 16'hD5D8, 16'hD619, 16'hE65A, 16'hE65A, 16'hDDD9, 16'h7A8B, 16'hA492, 16'hD619, 16'hC597, 16'hACD4, 16'hB555, 16'hC5D7, 16'hCE18,
        16'hC5D7, 16'hA492, 16'h9C51, 16'hA492, 16'h6249, 16'h72CB, 16'hB515, 16'hB555, 16'hCDD7, 16'h7B4D, 16'h730C, 16'h8B8E, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDE, 16'hCDD7, 16'h830B, 16'h6987, 16'hC556, 16'hE69B, 16'hEF1C, 16'hEF1D, 16'hEF1D, 16'hE71C, 16'hE6DB, 16'hE69A, 16'hA38E, 16'hC555, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF1E, 16'hFF5F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hD413, 16'hE5D8, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hF75D, 16'hFFDF, 16'hEEDC, 16'hEE5B, 16'hF69C, 16'hDD98, 16'hCD57, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hF69C, 16'hEE9C, 16'hF69C, 16'hAB4F, 16'hD557, 16'hFF1E, 16'hE558, 16'hE5D9, 16'hF69C, 16'hF69C, 16'hF6DD, 16'hE598, 16'hDDD8, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF69C, 16'hF69C, 16'hE5D9, 16'hE619, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hE619, 16'hBC53, 16'hE619, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B,
        16'hEE5B, 16'h8B0C, 16'h9B8F, 16'hE61A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hDDD8, 16'hBC94, 16'hDE19, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hE69B, 16'hE65A, 16'hB412, 16'h82CC, 16'hE619, 16'hE65B, 16'hE65A, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE1A, 16'hE65A, 16'hD5D9, 16'hD598, 16'hDE5A, 16'hE65A, 16'hE65A, 16'h9BD0, 16'h7B0C, 16'hCDD8, 16'hC5D8, 16'h7B4E, 16'h72CC, 16'h834E, 16'h8BCF, 16'h9C52, 16'h834E, 16'h3000, 16'h7B4D, 16'h8B8E, 16'h9C51, 16'hACD4, 16'hB515, 16'hCDD8, 16'h9C92, 16'h49C7, 16'h938F, 16'hACD4, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9B, 16'h82CB, 16'hDE59, 16'hE6DC, 16'hE6DB, 16'hD65A, 16'hD659, 16'hD659, 16'hD699, 16'hCD56, 16'h92CB, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5F, 16'hFF1E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF6DC, 16'hD3D2, 16'hF6DC, 16'hFFDF, 16'hFF9F, 16'hEE9B, 16'hEE9B, 16'hEEDC, 16'hEE5B, 16'hEE9B,
        16'hEE9B, 16'hD557, 16'hDD98, 16'hF69C, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hF6DC, 16'hEE1A, 16'h9A8C, 16'hEE1A, 16'hFF1D, 16'hE557, 16'hDD98, 16'hF69C, 16'hF69C, 16'hF6DD, 16'hDD98, 16'hDD98, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF69C, 16'hF69C, 16'hF69B, 16'hE5D9, 16'hE5D9, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE61A, 16'hC453, 16'hDD98, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hE65A, 16'hE61A, 16'hE61A, 16'hEE5A, 16'hA38F, 16'h7A4A, 16'hDDD9, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE65A, 16'hE61A, 16'hE65A, 16'hE61A, 16'hE61A, 16'hE65A, 16'hE619, 16'hBCD4, 16'hD598, 16'hEE9B, 16'hE69B, 16'hE65B, 16'hE69B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE69B, 16'hE65A, 16'hC4D4, 16'h79C9, 16'hCD97, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE1A, 16'hDE1A, 16'hDE1A, 16'hDE5A, 16'hDE19, 16'hDDD9, 16'hDE19, 16'hDE19,
        16'hCD97, 16'hDE5A, 16'hDE5A, 16'hE65A, 16'hC4D5, 16'h5986, 16'hA493, 16'hCE18, 16'hB514, 16'h8BCF, 16'hBD15, 16'hACD3, 16'hA492, 16'h9C51, 16'h9410, 16'hBD55, 16'hB515, 16'hA493, 16'hA492, 16'hACD4, 16'hCDD7, 16'hBD55, 16'h30C3, 16'h9C10, 16'h93CF, 16'hDE9B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC596, 16'hBD14, 16'hFF9E, 16'hE69B, 16'hD659, 16'hD659, 16'hD659, 16'hCE59, 16'hDE9A, 16'hA34D, 16'hDE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF1E, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hEE1A, 16'hD454, 16'hFF5E, 16'hFFDF, 16'hEEDC, 16'hE65B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hEE9C, 16'hE65A, 16'hCD16, 16'hE61A, 16'hF69C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hF6DC, 16'hDD98, 16'h9A8C, 16'hF69C, 16'hF6DD, 16'hDD57, 16'hDD97, 16'hEE9C, 16'hF69C, 16'hF6DC, 16'hDD98, 16'hDD98, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF69C, 16'hF69C, 16'hF69C, 16'hF69C, 16'hEE9B, 16'hEE9B, 16'hDDD9, 16'hDDD8, 16'hF69C, 16'hEE9B, 16'hEE9B,
        16'hEE9B, 16'hEE9B, 16'hEE5A, 16'hC453, 16'hD556, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hE61A, 16'hDDD9, 16'hDDD9, 16'hDDD8, 16'hEE1A, 16'hB410, 16'h4800, 16'hCD57, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE61A, 16'hE61A, 16'hBCD4, 16'hCD56, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hCD16, 16'h7A09, 16'hB4D4, 16'hE65A, 16'hE61A, 16'hE65A, 16'hDE1A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD9, 16'hD5D9, 16'hCD97, 16'hD5D8, 16'hCD97, 16'hD619, 16'hDE5A, 16'hDE5A, 16'hD598, 16'h7A8B, 16'h5186, 16'h7B4D, 16'hA492, 16'h6249, 16'hACD4, 16'hCDD8, 16'hCDD7, 16'hCDD7, 16'hC596, 16'hC596, 16'hBD55, 16'hA492, 16'h9C52, 16'hA493, 16'hC596, 16'hD5D8, 16'h7B4D, 16'h5208, 16'hB4D3, 16'h9C11, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA451, 16'hEEDB, 16'hCE18, 16'hACD3, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hC515, 16'hAC10, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5F, 16'hFEDD, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFF1E, 16'hFEDD, 16'hDD16, 16'hD4D5, 16'hFFDF, 16'hF75D, 16'hEE5A, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hE619, 16'hCD16, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hCCD5, 16'hA34F, 16'hFEDD, 16'hF6DC, 16'hD516, 16'hDD97, 16'hEE9B, 16'hEE9C, 16'hF69C, 16'hDD97, 16'hD557, 16'hF69C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF69C, 16'hF69C, 16'hF69C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hDDD8, 16'hDD98, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hC494, 16'hC4D4, 16'hEE5B, 16'hE65A, 16'hE65A, 16'hDE19, 16'hDDD8, 16'hD598, 16'hD597, 16'hDDD9, 16'hB411, 16'h2800, 16'hB493, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE619, 16'hC4D5, 16'hC515, 16'hDE19, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE61A, 16'hDE1A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hD597, 16'h8ACC, 16'h9BD0, 16'hE65A,
        16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD5D9, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD598, 16'hCD97, 16'hC557, 16'hCD97, 16'hD5D8, 16'hE65A, 16'hDE5A, 16'hDE19, 16'h938F, 16'h8B8E, 16'h938F, 16'h8B4E, 16'h8B8E, 16'hACD3, 16'hC597, 16'hC597, 16'hC596, 16'hC596, 16'hC556, 16'hC596, 16'hACD3, 16'h9C51, 16'h9C52, 16'hBD55, 16'hCDD8, 16'hAC93, 16'h000, 16'h93CF, 16'h9C10, 16'hC597, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hA410, 16'hC556, 16'h4040, 16'hACD3, 16'hDE5A, 16'hD659, 16'hCE19, 16'hDE59, 16'hA34D, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF1E, 16'hFF1E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hF6DD, 16'hF69C, 16'hCC13, 16'hDDD8, 16'hFFDF, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hDDD8, 16'hCD56, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF69C, 16'hBC12, 16'hABD0, 16'hFEDC, 16'hF69C, 16'hD516, 16'hD557, 16'hEE5B, 16'hEE9C, 16'hF69C, 16'hDD97, 16'hCD56, 16'hF69C, 16'hF69C, 16'hF69C, 16'hF69C, 16'hF69C, 16'hF69C, 16'hF69C, 16'hF69C, 16'hF69B, 16'hEE5B,
        16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5A, 16'hDD98, 16'hD557, 16'hEE5B, 16'hEE9B, 16'hEE5B, 16'hE65A, 16'hE65A, 16'hEE5A, 16'hC4D5, 16'hBC53, 16'hE619, 16'hE61A, 16'hE619, 16'hDDD8, 16'hD597, 16'hD597, 16'hCD57, 16'hDD98, 16'hB411, 16'h6000, 16'h934D, 16'hDDD9, 16'hDDD9, 16'hDDD8, 16'hD598, 16'hDDD8, 16'hD5D8, 16'hDDD9, 16'hDE19, 16'hE619, 16'hE65A, 16'hCD56, 16'hBCD4, 16'hD5D8, 16'hE65A, 16'hE61A, 16'hDE19, 16'hDDD9, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE61A, 16'hDD98, 16'hA34F, 16'h8B0C, 16'hDE19, 16'hDE19, 16'hD619, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hCD97, 16'hCD97, 16'hCD97, 16'hD5D8, 16'hCD97, 16'hCD97, 16'hC556, 16'hC556, 16'hCD97, 16'hDE1A, 16'hDE1A, 16'hE65A, 16'hAC52, 16'h8B4E, 16'hB4D4, 16'hAC52, 16'hAC51, 16'hC556, 16'hC597, 16'hC597, 16'hC597, 16'hC596, 16'hC596, 16'hC596, 16'hB515, 16'hA452, 16'h9C51, 16'hAD14, 16'hC5D7, 16'hBD55, 16'h628A, 16'h4145, 16'hA451, 16'h93CF, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h4840, 16'h728A, 16'h7289, 16'hC596, 16'hDE9A, 16'hCDD8, 16'hD619, 16'hBCD4, 16'hB451, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5F, 16'hFEDD, 16'hFF5E, 16'hFFDF, 16'hFF5E, 16'hFF1E, 16'hF69C, 16'hF69C, 16'hEE1A, 16'hBB91, 16'hEE5A, 16'hF71D, 16'hEE5B, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hD597, 16'hD597, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF65B, 16'h9B0E, 16'hBC93, 16'hF6DC, 16'hEE9C, 16'hD516, 16'hD557, 16'hE61A, 16'hEE9B, 16'hEE9C, 16'hD557, 16'hCD15, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hE65A, 16'hE61A, 16'hE65A, 16'hE65A, 16'hEE5A, 16'hEE5A, 16'hE65A, 16'hE61A, 16'hDD98, 16'hD557, 16'hEE5A, 16'hEE9B, 16'hE65A, 16'hE619, 16'hDE19, 16'hE61A, 16'hCD15, 16'hB412, 16'hDDD9, 16'hDE19, 16'hDDD8, 16'hD598, 16'hD597, 16'hD597, 16'hCD57, 16'hD597, 16'hAC10, 16'h928A, 16'h8A8B, 16'hBC93, 16'hAC11, 16'h9B8F, 16'h934E, 16'h934E, 16'h9B8F, 16'h9B8F, 16'hAC51, 16'hBCD4, 16'hD597, 16'hCD16, 16'hBCD4, 16'hD597, 16'hDDD9, 16'hDDD9, 16'hD5D8,
        16'hD597, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hDE19, 16'hDDD8, 16'hABD1, 16'h7A4A, 16'hCD97, 16'hDE19, 16'hD5D8, 16'hD5D8, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD57, 16'hCD97, 16'hCD97, 16'hCD57, 16'hC556, 16'hC556, 16'hC556, 16'hDE19, 16'hDE19, 16'hDE5A, 16'hC516, 16'h7A8B, 16'hC516, 16'hA451, 16'h9BCF, 16'hAC93, 16'hC597, 16'hC597, 16'hC596, 16'hC596, 16'hC596, 16'hC596, 16'hBD56, 16'hA492, 16'h9C52, 16'hA492, 16'hC596, 16'hCDD7, 16'h8BCF, 16'h8B8E, 16'h9410, 16'h93CF, 16'hB4D4, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD96, 16'h838E, 16'hD618, 16'h8B8E, 16'hDE9A, 16'hCDD7, 16'h8B8E, 16'hC514, 16'hA34D, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF1E, 16'hFEDD, 16'hFF9F, 16'hFF9F, 16'hF69C, 16'hF69C, 16'hEE5B, 16'hF69C, 16'hE5D9, 16'hBBD1, 16'hEE5A, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hD556, 16'hDDD8, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hEE5A, 16'h81C9, 16'hC4D4, 16'hF6DC, 16'hEE9B, 16'hCCD5, 16'hD557, 16'hDE19, 16'hEE9B, 16'hEE9C,
        16'hD557, 16'hC4D4, 16'hEE5A, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hE61A, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hD557, 16'hCD16, 16'hE61A, 16'hEE5B, 16'hDE19, 16'hD5D8, 16'hD598, 16'hDDD8, 16'hCD16, 16'hB411, 16'hD597, 16'hDDD8, 16'hD597, 16'hCD57, 16'hCD56, 16'hCD57, 16'hCD56, 16'hD557, 16'hB451, 16'h8208, 16'h5986, 16'h4882, 16'h7208, 16'h7A4A, 16'h82CC, 16'h82CC, 16'h82CC, 16'h82CC, 16'h828B, 16'h7A8B, 16'h82CC, 16'h8B0D, 16'h9B8F, 16'hC515, 16'hD5D8, 16'hD5D8, 16'hCD97, 16'hCD56, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hDE19, 16'hDDD8, 16'hBC52, 16'h8A8B, 16'hC515, 16'hDE19, 16'hD5D8, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hC556, 16'hCD56, 16'hCD97, 16'hCD57, 16'hC556, 16'hC556, 16'hC556, 16'hD5D8, 16'hDE5A, 16'hDE5A, 16'hD5D8, 16'h7A8B, 16'hBD15, 16'hB4D3, 16'hA410, 16'h9C10, 16'hC556, 16'hC597, 16'hC597, 16'hC596, 16'hC596, 16'hC596, 16'hC556, 16'hACD4, 16'hA492,
        16'h9C52, 16'hB515, 16'hCDD7, 16'hA492, 16'h838E, 16'hCD97, 16'h8B8E, 16'h8B4D, 16'hDE5A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hEF5D, 16'hFFDF, 16'hC5D7, 16'h9C10, 16'hACD3, 16'h9B8F, 16'h9B0D, 16'hAB8E, 16'hBC52, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFEDD, 16'hFF1E, 16'hFF9F, 16'hEE9C, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hF69C, 16'hDD57, 16'hBC12, 16'hE619, 16'hE65B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hEE5B, 16'hCD56, 16'hDDD9, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hE5D9, 16'h6003, 16'hCD15, 16'hF6DC, 16'hEE5B, 16'hCCD5, 16'hD557, 16'hDDD8, 16'hEE5B, 16'hEE9C, 16'hDD97, 16'hC494, 16'hE619, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE5A, 16'hE61A, 16'hE5D9, 16'hDDD9, 16'hDDD9, 16'hE619, 16'hE619, 16'hE619, 16'hE61A, 16'hE61A, 16'hE619, 16'hD557, 16'hCD16, 16'hDE19, 16'hEE5A, 16'hDDD8, 16'hCD57, 16'hCD57, 16'hD597, 16'hCD16, 16'hABD1, 16'hCD56, 16'hD598, 16'hD597, 16'hCD57, 16'hCD57, 16'hCD56, 16'hCD56, 16'hD557, 16'hAC11, 16'h5001, 16'h69C8, 16'h51C7, 16'h8B4E, 16'h8B8F, 16'h8B4E,
        16'h8B0D, 16'h82CC, 16'h7A8B, 16'h7A4A, 16'h724A, 16'h7A8B, 16'h82CC, 16'h7209, 16'h82CC, 16'hA452, 16'hCD56, 16'hD598, 16'hCD97, 16'hCD57, 16'hCD97, 16'hCD97, 16'hCD57, 16'hCD57, 16'hCD57, 16'hD5D8, 16'hDDD8, 16'hBC52, 16'h828B, 16'hB492, 16'hD618, 16'hCDD7, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD57, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hCD97, 16'hDE19, 16'hDE19, 16'hDE19, 16'h934E, 16'hA452, 16'hCD97, 16'hA451, 16'h938F, 16'hB4D4, 16'hC597, 16'hC597, 16'hC597, 16'hC596, 16'hC596, 16'hC596, 16'hB4D4, 16'hA492, 16'h9C52, 16'hB514, 16'hC596, 16'hBD55, 16'h59C7, 16'hDE9A, 16'hC556, 16'h82CC, 16'h9C11, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h6A8A, 16'h5986, 16'hACD2, 16'hEE9A, 16'h9B4D, 16'h8987, 16'hE65A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF1E, 16'hFEDD, 16'hFF5F, 16'hF6DD, 16'hE65A, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hF69B, 16'hCCD5, 16'hBC93, 16'hE61A, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hE61A, 16'hCD16, 16'hDE19, 16'hEE5B, 16'hEE5B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65A,
        16'hE65A, 16'hEE5B, 16'hCD15, 16'h3800, 16'hD556, 16'hEE9C, 16'hE61A, 16'hC494, 16'hD557, 16'hDDD8, 16'hE619, 16'hEE9B, 16'hD597, 16'hBC53, 16'hDDD8, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hE61A, 16'hE619, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hE619, 16'hE619, 16'hDDD9, 16'hDDD8, 16'hD557, 16'hC4D5, 16'hDDD8, 16'hE61A, 16'hCD97, 16'hCD56, 16'hCD56, 16'hD557, 16'hCD16, 16'hABD1, 16'hCD15, 16'hD597, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD56, 16'hD597, 16'hAC10, 16'hA30D, 16'hE494, 16'h8ACC, 16'hD597, 16'hD5D8, 16'hD598, 16'hD598, 16'hCD57, 16'hBD15, 16'hBCD4, 16'hAC52, 16'h9BD0, 16'h934E, 16'h7A4A, 16'h7A8A, 16'h7A4A, 16'h82CC, 16'hAC51, 16'hCD56, 16'hCD97, 16'hC556, 16'hC556, 16'hC556, 16'hCD56, 16'hCD56, 16'hCD97, 16'hD598, 16'hB452, 16'h9B4E, 16'h9BD0, 16'hD5D8, 16'hCDD8, 16'hCDD7, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hC556, 16'hC556, 16'hC596, 16'hC596, 16'hC556, 16'hC556, 16'hC597, 16'hDE19, 16'hDE19, 16'hDE5A, 16'hAC52, 16'h8B8E,
        16'hDE19, 16'hBCD4, 16'h9B8F, 16'hA452, 16'hCD97, 16'hC596, 16'hC597, 16'hC596, 16'hC596, 16'hC596, 16'hBD55, 16'hA492, 16'hA492, 16'hACD3, 16'hBD96, 16'hCDD7, 16'h7B0C, 16'hB596, 16'hFF9E, 16'h9BD0, 16'h830C, 16'hBD95, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hB514, 16'hD5D7, 16'hFFDF, 16'hD597, 16'h3800, 16'hA410, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFEDD, 16'hFEDD, 16'hF71E, 16'hE65B, 16'hE65A, 16'hE65B, 16'hEE5B, 16'hEE9B, 16'hEE5A, 16'hBC52, 16'hC4D4, 16'hE65A, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hDE19, 16'hCD16, 16'hE61A, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hEE5B, 16'hA3D1, 16'h3800, 16'hD515, 16'hEE5B, 16'hDE19, 16'hC494, 16'hD557, 16'hD597, 16'hDDD8, 16'hEE5B, 16'hD597, 16'hBC93, 16'hD597, 16'hEE9B, 16'hEE5B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE619, 16'hDDD8, 16'hD598, 16'hD598, 16'hD598, 16'hD597, 16'hD598, 16'hDDD9, 16'hDDD8, 16'hD597, 16'hD597, 16'hCD16, 16'hC4D5, 16'hD597, 16'hDDD8, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hABD1, 16'hC4D5, 16'hD597, 16'hCD57,
        16'hCD57, 16'hCD57, 16'hCD56, 16'hCD56, 16'hD597, 16'hA3D0, 16'hAB0D, 16'hED16, 16'h9ACC, 16'hAC52, 16'hDDD8, 16'hD598, 16'hD598, 16'hD598, 16'hD598, 16'hD5D8, 16'hD5D8, 16'hD597, 16'hD597, 16'hB452, 16'hA3D1, 16'hAC52, 16'h934E, 16'h724A, 16'h7ACC, 16'hB493, 16'hCD56, 16'hCD56, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hD597, 16'hB452, 16'hABD0, 16'h934E, 16'hD598, 16'hD5D8, 16'hCDD7, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD57, 16'hC556, 16'hC596, 16'hC596, 16'hC556, 16'hC556, 16'hC556, 16'hD619, 16'hDE59, 16'hE65A, 16'hC515, 16'h7ACC, 16'hD619, 16'hCD97, 16'hA411, 16'h93D0, 16'hC597, 16'hC597, 16'hC596, 16'hC597, 16'hC596, 16'hC596, 16'hC596, 16'hACD3, 16'hA492, 16'hA4D3, 16'hB514, 16'hCDD7, 16'hA452, 16'h7B4D, 16'hFFDF, 16'hE6DB, 16'h830C, 16'h7ACC, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hFF9E, 16'hEE9B, 16'h92CB, 16'h6000, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hFE9D, 16'hFEDD, 16'hEE5B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65B, 16'hEE9B, 16'hE619, 16'hB411, 16'hCD56, 16'hE65A, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B,
        16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hD598, 16'hCD56, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE61A, 16'hE65A, 16'hE5D9, 16'h7A4A, 16'h6145, 16'hCD15, 16'hE61A, 16'hDDD9, 16'hC494, 16'hD557, 16'hD597, 16'hD597, 16'hDDD9, 16'hD557, 16'hBC93, 16'hCD56, 16'hE61A, 16'hE61A, 16'hE65A, 16'hE65A, 16'hE61A, 16'hDDD8, 16'hD597, 16'hD597, 16'hD557, 16'hD557, 16'hD557, 16'hD597, 16'hDDD8, 16'hD598, 16'hCD56, 16'hCD56, 16'hCD16, 16'hC4D5, 16'hCD57, 16'hD597, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hD556, 16'hB3D1, 16'hBC93, 16'hD597, 16'hCD56, 16'hCD57, 16'hCD57, 16'hCD56, 16'hCD56, 16'hD597, 16'hA3CF, 16'hB34E, 16'hECD6, 16'hC3D1, 16'h934D, 16'hD5D8, 16'hD598, 16'hD597, 16'hCD97, 16'hD597, 16'hCD97, 16'hCD97, 16'hCD57, 16'hD598, 16'hC4D4, 16'hB452, 16'hD5D8, 16'hCD56, 16'hBCD5, 16'hA411, 16'h8B0D, 16'h938E, 16'hBCD4, 16'hCD56, 16'hC516, 16'hC516, 16'hC556, 16'hCD97, 16'hB452, 16'hB411, 16'h8B0D, 16'hCD97, 16'hD5D8, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97,
        16'hCD97, 16'hCD56, 16'hC556, 16'hCD96, 16'hC556, 16'hC557, 16'hC556, 16'hD5D8, 16'hDE59, 16'hDE5A, 16'hCD97, 16'h724A, 16'hCD97, 16'hDE19, 16'hB493, 16'h938E, 16'hBD15, 16'hCD97, 16'hC596, 16'hC596, 16'hC597, 16'hC597, 16'hC596, 16'hACD4, 16'hA493, 16'hA492, 16'hACD4, 16'hC597, 16'hB515, 16'h5A08, 16'hE71C, 16'hFFDF, 16'hD618, 16'h6A09, 16'h93D0, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'hE6DB, 16'hEF1C, 16'hCD15, 16'hC452, 16'hC4D4, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFEDD, 16'hFEDD, 16'hF69C, 16'hE61A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hDDD8, 16'hB3D1, 16'hCD56, 16'hE65A, 16'hE65B, 16'hE65B, 16'hE65A, 16'hE65B, 16'hE65A, 16'hE65B, 16'hE65B, 16'hCD57, 16'hD557, 16'hE65A, 16'hE61A, 16'hE61A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE61A, 16'hCD56, 16'h6145, 16'h7A09, 16'hCD15, 16'hDDD9, 16'hDDD8, 16'hC4D4, 16'hD556, 16'hD557, 16'hD597, 16'hD597, 16'hD557, 16'hC493, 16'hCD15, 16'hDDD8, 16'hDDD8, 16'hE65A, 16'hE61A, 16'hE619, 16'hDD98, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hCD57, 16'hCD57, 16'hD597, 16'hCD57, 16'hCD16, 16'hCD16, 16'hC515,
        16'hC4D5, 16'hCD56, 16'hD597, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hD557, 16'hB412, 16'hB411, 16'hD597, 16'hCD57, 16'hCD57, 16'hCD56, 16'hCD56, 16'hC556, 16'hD597, 16'hA38F, 16'hBBD1, 16'hED17, 16'hE494, 16'h928B, 16'hCD15, 16'hD598, 16'hD597, 16'hCD97, 16'hCD97, 16'hCD97, 16'hD597, 16'hCD97, 16'hD598, 16'hCD15, 16'hA38F, 16'hCD56, 16'hCD97, 16'hCD57, 16'hCD57, 16'hCD56, 16'hBC93, 16'hA3D0, 16'hB493, 16'hC515, 16'hC556, 16'hC556, 16'hCD57, 16'hB492, 16'hB411, 16'h934D, 16'hBD15, 16'hD5D9, 16'hD5D8, 16'hD5D8, 16'hCD98, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD57, 16'hCD96, 16'hCD97, 16'hC557, 16'hC556, 16'hC556, 16'hCDD7, 16'hDE19, 16'hDE5A, 16'hDE19, 16'h830D, 16'hB514, 16'hDE5A, 16'hC556, 16'h938E, 16'hB4D4, 16'hCD97, 16'hC597, 16'hC596, 16'hC596, 16'hC596, 16'hCD97, 16'hB515, 16'hA493, 16'hA492, 16'hACD3, 16'hBD56, 16'hC597, 16'h6208, 16'hC596, 16'hFFDF, 16'hFFDF, 16'hB555, 16'h5004, 16'hC596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'hDE59, 16'hF6DB, 16'hC514, 16'hEEDB, 16'hA34E, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFF5E, 16'hFFDF, 16'hFF5E, 16'hFEDC, 16'hFE9D, 16'hE61A, 16'hE61A, 16'hE65A,
        16'hE65A, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hD557, 16'hABD1, 16'hCD56, 16'hDE19, 16'hE65B, 16'hE65A, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE61A, 16'hCD56, 16'hD597, 16'hE61A, 16'hE61A, 16'hDE19, 16'hDDD9, 16'hDDD9, 16'hDE19, 16'hDDD9, 16'hE61A, 16'hAC12, 16'h6946, 16'h824A, 16'hCD15, 16'hD598, 16'hD597, 16'hC4D4, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD57, 16'hD557, 16'hC4D4, 16'hC4D4, 16'hD597, 16'hD557, 16'hDDD8, 16'hE619, 16'hD598, 16'hD597, 16'hD597, 16'hCD57, 16'hD597, 16'hCD56, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD56, 16'hC515, 16'hCD16, 16'hC515, 16'hC4D5, 16'hCD56, 16'hD557, 16'hCD56, 16'hCD16, 16'hCD56, 16'hCD56, 16'hD557, 16'hB412, 16'hABD1, 16'hD597, 16'hD597, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD56, 16'hD597, 16'h9B4E, 16'hC453, 16'hED17, 16'hECD6, 16'hAB4E, 16'hAC51, 16'hDDD8, 16'hD597, 16'hCD97, 16'hCD97, 16'hCD57, 16'hD597, 16'hCD97, 16'hD597, 16'hD556, 16'hA38F, 16'hCD56, 16'hCD97, 16'hCD56, 16'hC556, 16'hC556, 16'hCD97, 16'hCD56, 16'hC515, 16'hB494, 16'hBD15, 16'hC556,
        16'hCD57, 16'hB493, 16'hAC11, 16'h9B4E, 16'hBCD4, 16'hDE19, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hCD98, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD57, 16'hCD97, 16'hCD97, 16'hDE19, 16'hDE5A, 16'hDE5A, 16'h9BD0, 16'hAC52, 16'hDE19, 16'hD5D8, 16'h9BD0, 16'hA411, 16'hCD97, 16'hC597, 16'hC597, 16'hC596, 16'hC596, 16'hCD97, 16'hBD55, 16'hA493, 16'hA492, 16'hA493, 16'hB514, 16'hC5D7, 16'h8BCF, 16'h8BCF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'h93CF, 16'h6A49, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD618, 16'hD5D7, 16'hEEDB, 16'hBC93, 16'hFF5E, 16'hCD56, 16'hB493, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF6DC, 16'hFF9E, 16'hFFDF, 16'hFF1D, 16'hFE9C, 16'hF69C, 16'hDE19, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE65A, 16'hE65A, 16'hEE5B, 16'hCD16, 16'hB452, 16'hD597, 16'hDE19, 16'hE65A, 16'hDE19, 16'hE61A, 16'hDE19, 16'hDE19, 16'hE61A, 16'hDE19, 16'hCD15, 16'hD597, 16'hDE19, 16'hDDD9, 16'hDDD9, 16'hDE19, 16'hE619, 16'hDDD8, 16'hD597, 16'hD597, 16'h7A8B, 16'hA30D, 16'h828B, 16'hC515, 16'hD597, 16'hCD56, 16'hC4D4, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD56, 16'hCD57, 16'hC4D5, 16'hC4D4, 16'hCD16, 16'hCD16, 16'hCD56, 16'hD597, 16'hD597,
        16'hD597, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD56, 16'hCD57, 16'hCD56, 16'hC515, 16'hCD16, 16'hC515, 16'hC4D5, 16'hCD56, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD16, 16'hCD56, 16'hD557, 16'hBC53, 16'hAB90, 16'hD557, 16'hD597, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hD557, 16'h930D, 16'hD494, 16'hED58, 16'hE495, 16'hCC13, 16'h930D, 16'hDDD8, 16'hD597, 16'hCD57, 16'hD597, 16'hCD97, 16'hD597, 16'hD597, 16'hD597, 16'hD557, 16'h9B4F, 16'hC515, 16'hCD97, 16'hCD56, 16'hCD56, 16'hC556, 16'hC556, 16'hCD56, 16'hCD56, 16'hC556, 16'hC515, 16'hC556, 16'hCD56, 16'hBC93, 16'hABD0, 16'hABD0, 16'hB452, 16'hDE19, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD598, 16'hD597, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hD619, 16'hDE59, 16'hE65A, 16'hB493, 16'h8B4E, 16'hDE19, 16'hDE19, 16'hAC93, 16'h8B4E, 16'hC597, 16'hC597, 16'hC597, 16'hC597, 16'hC596, 16'hCDD7, 16'hC596, 16'hA492, 16'hA492, 16'hA492, 16'hACD4, 16'hC596, 16'hACD3, 16'h5A08, 16'hEF1D,
        16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h5986, 16'hA492, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCDD7, 16'hD5D7, 16'hEE5A, 16'hB452, 16'hF71D, 16'hFF5E, 16'hA38F, 16'hF75D, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFF1D, 16'hEE9B, 16'hFFDF, 16'hFF9F, 16'hFEDD, 16'hFE9D, 16'hE61A, 16'hD5D8, 16'hE61A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE61A, 16'hE65A, 16'hC4D4, 16'hBC53, 16'hD597, 16'hDDD9, 16'hDDD9, 16'hD5D8, 16'hD5D8, 16'hD598, 16'hDDD8, 16'hDDD9, 16'hD5D8, 16'hC515, 16'hDD97, 16'hDE19, 16'hDE19, 16'hDDD8, 16'hC515, 16'hAC11, 16'h9B8F, 16'h934E, 16'h82CC, 16'h3882, 16'hAB8F, 16'h7A49, 16'hC515, 16'hD597, 16'hCD56, 16'hC4D4, 16'hCD16, 16'hCD16, 16'hCD16, 16'hCD56, 16'hCD56, 16'hCD15, 16'hC4D4, 16'hC515, 16'hCD16, 16'hCD56, 16'hCD56, 16'hCD57, 16'hD597, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD57, 16'hCD56, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hCD56, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hD597, 16'hBC94, 16'hAB4F, 16'hCD56, 16'hCD97, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hD597, 16'h9B0C, 16'hDCD5, 16'hF599, 16'hE4D5, 16'hED16, 16'h928B, 16'hCD15, 16'hD598, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hDD97,
        16'h9B4E, 16'hC4D4, 16'hCD97, 16'hCD56, 16'hCD56, 16'hC556, 16'hCD56, 16'hCD56, 16'hC556, 16'hCD56, 16'hC556, 16'hC516, 16'hC556, 16'hBCD4, 16'hA34E, 16'hAC11, 16'h9BCF, 16'hDE19, 16'hD5D9, 16'hD5D9, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD598, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hD5D8, 16'hDE59, 16'hE65A, 16'hC515, 16'h830D, 16'hD5D8, 16'hDE19, 16'hC556, 16'h82CC, 16'hBD15, 16'hC597, 16'hC597, 16'hC596, 16'hC596, 16'hC597, 16'hC597, 16'hACD3, 16'hA492, 16'hA492, 16'hACD3, 16'hBD55, 16'hBD56, 16'h5A08, 16'hCE19, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE18, 16'h3800, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD97, 16'hDE18, 16'hE619, 16'hB411, 16'hEF1C, 16'hFFDF, 16'hC515, 16'hCDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE1A, 16'hF6DC, 16'hFFDF, 16'hFF5E, 16'hFE9C, 16'hFE9C, 16'hDDD9, 16'hD598, 16'hDDD9, 16'hD598, 16'hD5D8, 16'hDDD9, 16'hD5D8, 16'hDE19, 16'hBC93, 16'hBC93, 16'hD597, 16'hD597, 16'hCD56, 16'hCD56, 16'hCD97, 16'hCD56, 16'hCD57, 16'hD597, 16'hCD97, 16'hC515, 16'hDDD8, 16'hDDD8, 16'hBD15, 16'h934F, 16'h828B, 16'h828B, 16'h7A4B, 16'h7209, 16'h5146, 16'h4145, 16'h8ACC, 16'h69C7, 16'hC515, 16'hCD97, 16'hCD56, 16'hC4D4,
        16'hCD15, 16'hC515, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD16, 16'hC4D4, 16'hC515, 16'hC516, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD57, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hCD56, 16'hCD97, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hD597, 16'hC4D4, 16'hA30E, 16'hC515, 16'hD597, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD56, 16'hD556, 16'h9A8B, 16'hDD16, 16'hFE1B, 16'hE557, 16'hF557, 16'hBBD1, 16'hAC11, 16'hDDD8, 16'hD598, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hDD97, 16'h9B0D, 16'hBC93, 16'hCD97, 16'hCD96, 16'hCD96, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hC555, 16'hC556, 16'hC556, 16'hC4D4, 16'h9B4E, 16'hB452, 16'hA3D0, 16'hDDD9, 16'hD619, 16'hDE19, 16'hDDD9, 16'hD5D9, 16'hD5D9, 16'hD5D8, 16'hD5D8, 16'hD598, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hD5D8, 16'hDE59, 16'hE65A, 16'hCD97, 16'h830C, 16'hCD97, 16'hDE59, 16'hD618, 16'h8B0D, 16'hAC93, 16'hCDD7, 16'hCD97,
        16'hCD97, 16'hC597, 16'hC597, 16'hC597, 16'hACD4, 16'hA492, 16'hA493, 16'hA492, 16'hACD4, 16'hC596, 16'h7B0C, 16'h9C51, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hACD3, 16'h6208, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFF9E, 16'hCD56, 16'hE619, 16'hDDD8, 16'hB492, 16'hF75D, 16'hFFDF, 16'hF71C, 16'hB452, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hE599, 16'hFF9E, 16'hFFDF, 16'hFEDD, 16'hF69C, 16'hF69B, 16'hCD97, 16'hD598, 16'hCD97, 16'hC556, 16'hCD97, 16'hCD97, 16'hCD57, 16'hD5D8, 16'hBC93, 16'hBCD4, 16'hCD97, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD97, 16'hCD16, 16'hCD16, 16'hC515, 16'h9B8F, 16'h828B, 16'h828B, 16'h828B, 16'h82CC, 16'h9B8F, 16'hB493, 16'h6249, 16'hB411, 16'hF557, 16'h7A09, 16'hC515, 16'hD557, 16'hCD16, 16'hBC93, 16'hCD15, 16'hC516, 16'hCD16, 16'hCD56, 16'hCD56, 16'hCD56, 16'hBC94, 16'hCD15, 16'hCD16, 16'hC516, 16'hC515, 16'hCD56, 16'hCD57, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC515, 16'hC515, 16'hC515, 16'hC515, 16'hCD56, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD15, 16'hA2CE, 16'hC494, 16'hD597, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD57, 16'hCD56, 16'h924A, 16'hE557, 16'hFE9C,
        16'hF65B, 16'hED17, 16'hE516, 16'h930C, 16'hDD98, 16'hD598, 16'hD597, 16'hD598, 16'hD597, 16'hD597, 16'hD597, 16'hDD98, 16'h9B4E, 16'hA3D1, 16'hD597, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC556, 16'hCD56, 16'hC556, 16'hCD56, 16'hC516, 16'hCD56, 16'hC515, 16'h9B0D, 16'hBC53, 16'h934E, 16'hDDD9, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD5D9, 16'hDDD9, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD98, 16'hDE59, 16'hE69A, 16'hDE19, 16'h8B0E, 16'hC556, 16'hDE59, 16'hDE19, 16'hAC12, 16'h938F, 16'hCDD7, 16'hCD97, 16'hC597, 16'hC597, 16'hC597, 16'hCDD7, 16'hB514, 16'hA492, 16'hA493, 16'hA492, 16'hACD3, 16'hBD55, 16'h9C51, 16'h6249, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h72CB, 16'h9BD0, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hCD55, 16'hEE5A, 16'hD597, 16'hBC93, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hC514, 16'hDE59, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hE5D9, 16'hEE1A, 16'hFFDF, 16'hFF5E, 16'hF69C, 16'hF69C, 16'hE619, 16'hC556, 16'hCD57, 16'hCD56, 16'hC556, 16'hC556, 16'hCD56, 16'hCD56, 16'hD597, 16'hB452, 16'hC4D4, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC556, 16'hCD56, 16'hCD57, 16'hCD15, 16'hA390, 16'h8ACC, 16'h7A8B, 16'h7A8B, 16'h82CC,
        16'hAC52, 16'hC515, 16'hCD97, 16'hD597, 16'h7A4A, 16'hD4D4, 16'hED16, 16'h7A09, 16'hC4D5, 16'hD598, 16'hCD16, 16'hB412, 16'hCD16, 16'hC515, 16'hC515, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC494, 16'hCD15, 16'hCD16, 16'hC515, 16'hCD16, 16'hCD16, 16'hCD56, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD57, 16'hCD57, 16'hCD56, 16'hC516, 16'hC515, 16'hC515, 16'hC515, 16'hCD56, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hD557, 16'hCD16, 16'h924C, 16'hC453, 16'hD597, 16'hD557, 16'hCD57, 16'hCD56, 16'hD597, 16'hCD16, 16'h928B, 16'hED57, 16'hFE9C, 16'hFF1E, 16'hED57, 16'hF558, 16'hA30E, 16'hCCD4, 16'hDDD8, 16'hDD98, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hD598, 16'hE5D8, 16'h9B4E, 16'h828B, 16'hD556, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC515, 16'h930D, 16'hC493, 16'h930D, 16'hDDD8, 16'hDE5A, 16'hDE5A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hCD97, 16'hD597, 16'hD598,
        16'hCD98, 16'hDE19, 16'hDE5A, 16'hDE1A, 16'h934F, 16'hB493, 16'hDE59, 16'hDE19, 16'hC515, 16'h7A8B, 16'hC597, 16'hCDD7, 16'hC597, 16'hC597, 16'hC597, 16'hCDD7, 16'hBD55, 16'hA492, 16'hA492, 16'hA492, 16'hA493, 16'hB514, 16'hB514, 16'h4985, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h3000, 16'hBD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'hCD15, 16'hEE5A, 16'hD516, 16'hBD14, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hB492, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hEE9C, 16'hDD57, 16'hEEDC, 16'hFFDF, 16'hFF1D, 16'hF69B, 16'hF69B, 16'hD598, 16'hC556, 16'hCD56, 16'hCD56, 16'hC556, 16'hC556, 16'hC556, 16'hC556, 16'hD597, 16'hB452, 16'hC515, 16'hCD97, 16'hCD56, 16'hCD56, 16'hC556, 16'hC556, 16'hCD56, 16'hCD57, 16'hC515, 16'h9B4E, 16'h828B, 16'h828C, 16'h82CC, 16'hAC52, 16'hCD56, 16'hD597, 16'hCD97, 16'hD5D7, 16'hBC93, 16'h8209, 16'hED16, 16'hED58, 16'h8B0D, 16'hC4D4, 16'hDD98, 16'hCD16, 16'hAC11, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD57, 16'hC494, 16'hCD15, 16'hCD16, 16'hCD16, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD57, 16'hCD56, 16'hCD57, 16'hCD57, 16'hCD56, 16'hC516, 16'hCD16, 16'hC516, 16'hCD16, 16'hD597, 16'hD597, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD16, 16'hD557,
        16'hD556, 16'h924B, 16'hBC11, 16'hDD97, 16'hD597, 16'hD597, 16'hD557, 16'hD597, 16'hCCD5, 16'hA2CC, 16'hF598, 16'hF6DC, 16'hFF9F, 16'hF5D9, 16'hF558, 16'hCC53, 16'hABD0, 16'hE5D9, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hE5D8, 16'hB3D0, 16'h7041, 16'hC493, 16'hD597, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD57, 16'hCD16, 16'h9B0D, 16'hC453, 16'h8B0D, 16'hD597, 16'hDE5A, 16'hDE5A, 16'hDE5A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD5D8, 16'hD5D8, 16'hCD98, 16'hD5D8, 16'hD5D8, 16'hD598, 16'hDE19, 16'hDE5A, 16'hE65A, 16'hA3D1, 16'hAC52, 16'hDE5A, 16'hD619, 16'hD5D8, 16'h7A8B, 16'hBD15, 16'hCDD8, 16'hCDD7, 16'hC597, 16'hC596, 16'hC597, 16'hBD56, 16'hA492, 16'hA492, 16'hA492, 16'hA492, 16'hACD3, 16'hBD55, 16'h628A, 16'h9C92, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD96, 16'h2800, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65A, 16'hCCD4, 16'hF69B, 16'hCD15, 16'hC555, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD96, 16'hDE5A, 16'hFFDF, 16'hFF5E, 16'hFFDF, 16'hFF5E, 16'hE5D9, 16'hDD97, 16'hF71D, 16'hFFDF, 16'hF6DC, 16'hEE5B, 16'hEE5A, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC556, 16'hCD56, 16'hCD56, 16'hCD57, 16'hCD97, 16'hB452, 16'hC515, 16'hCD57, 16'hCD56,
        16'hCD56, 16'hC556, 16'hCD56, 16'hCD57, 16'hC515, 16'h930D, 16'h6A09, 16'h8ACC, 16'hAC11, 16'hCD16, 16'hD598, 16'hCD97, 16'hCD97, 16'hCD97, 16'hD598, 16'hA3D0, 16'hAB0E, 16'hED17, 16'hF61A, 16'hA411, 16'hBC93, 16'hDD98, 16'hCD16, 16'h9B0E, 16'hCD15, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD57, 16'hC4D4, 16'hC4D4, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD57, 16'hCD56, 16'hCD57, 16'hD597, 16'hCD57, 16'hCD57, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hD597, 16'hD597, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hD597, 16'hD556, 16'h920A, 16'hB3D0, 16'hDD98, 16'hD597, 16'hD597, 16'hD597, 16'hDDD8, 16'hC4D4, 16'hAACD, 16'hF5D9, 16'hFEDD, 16'hFF9F, 16'hFE9C, 16'hF558, 16'hE517, 16'h9ACC, 16'hDD97, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hE5D9, 16'hB410, 16'h9A4A, 16'h9B0D, 16'hDD97, 16'hD597, 16'hCD97, 16'hCD57, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'h92CC, 16'hC452, 16'h934D, 16'hCD97, 16'hE65A, 16'hDE5A,
        16'hE65A, 16'hDE5A, 16'hDE5A, 16'hDE1A, 16'hDE19, 16'hDE1A, 16'hDE1A, 16'hD5D9, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hDE19, 16'hDE5A, 16'hE65A, 16'hB493, 16'h93D0, 16'hDE19, 16'hDE19, 16'hDE19, 16'h8B0E, 16'hAC92, 16'hCDD8, 16'hC597, 16'hC596, 16'hC596, 16'hC596, 16'hC596, 16'hACD3, 16'hA492, 16'hA492, 16'hA492, 16'hA492, 16'hB555, 16'h8B8F, 16'h6ACA, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h93D0, 16'h728A, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD5D8, 16'hCD16, 16'hF69B, 16'hC4D4, 16'hCDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hBC93, 16'hFFDF, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hEE5B, 16'hD557, 16'hDDD8, 16'hFF5E, 16'hFF5E, 16'hEE9B, 16'hEE9B, 16'hE619, 16'hCD56, 16'hCD57, 16'hCD57, 16'hCD97, 16'hCD56, 16'hCD57, 16'hCD56, 16'hCD97, 16'hCD97, 16'hAC12, 16'hC515, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD57, 16'hC515, 16'h8ACC, 16'h824A, 16'h8B0D, 16'hBCD5, 16'hD5D8, 16'hD597, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hD597, 16'h828C, 16'hCC12, 16'hED16, 16'hFEDD, 16'hAC93, 16'hAC11, 16'hDDD8, 16'hD556, 16'h7A09, 16'hC4D4, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD56, 16'hD597, 16'hC4D5, 16'hC493, 16'hD557, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD57, 16'hD597, 16'hD597, 16'hD597, 16'hD597,
        16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hD557, 16'hDD98, 16'hD597, 16'hCD56, 16'hCD56, 16'hD556, 16'hD557, 16'hD597, 16'hDD57, 16'h920A, 16'hA34E, 16'hDDD8, 16'hD597, 16'hDDD8, 16'hDD97, 16'hE5D9, 16'hBC53, 16'hB34F, 16'hFDD9, 16'hFF1E, 16'hFF9F, 16'hFF5E, 16'hED99, 16'hF599, 16'hB3D0, 16'hC493, 16'hE5D9, 16'hDDD8, 16'hE5D8, 16'hE5D9, 16'hDDD8, 16'hEDD9, 16'hB3D0, 16'hC391, 16'h9A8C, 16'hBC93, 16'hDD98, 16'hD597, 16'hD597, 16'hCD97, 16'hD597, 16'hCD57, 16'hCD57, 16'hCD97, 16'hCD97, 16'hD597, 16'h92CC, 16'hBC11, 16'h9B4E, 16'hCD56, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE1A, 16'hDE5A, 16'hDE19, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D9, 16'hDE5A, 16'hE65B, 16'hC4D5, 16'h8B4D, 16'hDE19, 16'hDE19, 16'hDE5A, 16'hA452, 16'h93CF, 16'hCDD8, 16'hC597, 16'hC596, 16'hC597, 16'hC596, 16'hC596, 16'hBD55, 16'h9C52, 16'hA492, 16'hA493, 16'hA492, 16'hAD14, 16'hA492, 16'h2800, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D,
        16'h6208, 16'hA452, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD56, 16'hD557, 16'hEE5A, 16'hC493, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC4D4, 16'hE69B, 16'hFF9F, 16'hFF1E, 16'hFF5F, 16'hF69C, 16'hE5D9, 16'hD556, 16'hE61A, 16'hFF5F, 16'hF6DC, 16'hE65A, 16'hEE9B, 16'hDDD9, 16'hCD56,
        16'hCD97, 16'hCD97, 16'hCD97, 16'hCD57, 16'hCD57, 16'hCD97, 16'hD597, 16'hCD97, 16'hAC12, 16'hCD15, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hC515, 16'h82CC, 16'h82CC, 16'hBC94, 16'hBC94, 16'hCD57, 16'hD597, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD57, 16'hD597, 16'hCD15, 16'h81C9, 16'hE4D5, 16'hED57, 16'hFF5F, 16'hC516, 16'hA38F, 16'hDDD8, 16'hD556, 16'h6946, 16'hAC11, 16'hD597, 16'hD597, 16'hCD57, 16'hCD56, 16'hD598, 16'hCD16, 16'hB412, 16'hD557, 16'hCD56, 16'hCD16, 16'hCD56, 16'hCD56, 16'hCD57, 16'hCD57, 16'hCD57, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hCD56, 16'hCD57, 16'hD557, 16'hD597, 16'hDDD8, 16'hD597, 16'hD557, 16'hD557, 16'hD557, 16'hD557, 16'hD597, 16'hDD97, 16'h924B, 16'h928C, 16'hE5D8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hE619, 16'hABD0, 16'hCC11, 16'hFE1A, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hF69C, 16'hF598, 16'hE4D6, 16'hA30D, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hEDD9, 16'hAB90, 16'hCC12, 16'hCC12, 16'h930D, 16'hDDD8, 16'hD597, 16'hD597, 16'hD597,
        16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'h8A8C, 16'hC453, 16'h9B4E, 16'hCD56, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE1A, 16'hD5D9, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hDE5A, 16'hE69B, 16'hCD56, 16'h8B0D, 16'hDE19, 16'hDE19, 16'hDE5A, 16'hBD16, 16'h7ACC, 16'hCDD7, 16'hCDD7, 16'hC597, 16'hC597, 16'hC596, 16'hB555, 16'hBD56, 16'hA492, 16'hA492, 16'hA4D3, 16'hA4D3, 16'hA4D3, 16'hAD13, 16'h4144, 16'hA4D3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h3800, 16'hCD97, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hBD14, 16'hDDD8, 16'hE61A, 16'hC4D4, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hBCD3, 16'hFFDF, 16'hFF5E, 16'hFF5E, 16'hF6DC, 16'hEE5A, 16'hD598, 16'hD556, 16'hEE5B, 16'hFF5E, 16'hE65B, 16'hE65B, 16'hE65A, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hB452, 16'hCD56, 16'hCD57, 16'hC556, 16'hC556, 16'hCD56, 16'h9B8F, 16'h9B8F, 16'hC515, 16'hCD57, 16'hBC53, 16'hCD56, 16'hD598, 16'hCD97, 16'hD597, 16'hCD97, 16'hCD97, 16'hD598, 16'hB452, 16'h9A8C, 16'hED17, 16'hEDD9, 16'hFF9F, 16'hDE19, 16'h9B4E, 16'hDDD8, 16'hD556, 16'h824A, 16'h9B0D, 16'hD557, 16'hD597, 16'hCD97, 16'hD597, 16'hD598, 16'hD557, 16'hB3D0,
        16'hD557, 16'hD557, 16'hCD57, 16'hCD56, 16'hCD57, 16'hCD57, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hD557, 16'hD557, 16'hD597, 16'hDDD8, 16'hE5D9, 16'hDD98, 16'hD597, 16'hDD97, 16'hDD97, 16'hD597, 16'hDD98, 16'hDD97, 16'h9A8B, 16'h89C9, 16'hDD98, 16'hE619, 16'hDDD8, 16'hDDD9, 16'hE619, 16'hA30D, 16'hDC94, 16'hF65B, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hF5D9, 16'hF599, 16'hA30E, 16'hD516, 16'hEDD9, 16'hE5D8, 16'hE619, 16'hE5D9, 16'hEDD9, 16'hAB4E, 16'hD4D5, 16'hED16, 16'h9A8B, 16'hC4D4, 16'hE5D9, 16'hD598, 16'hD598, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'h92CC, 16'hC453, 16'hAB90, 16'hC556, 16'hE69B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE19, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D9, 16'hD5D8, 16'hDE5A, 16'hE69A, 16'hD597, 16'h830C, 16'hD597, 16'hDE19, 16'hDE19, 16'hD5D8, 16'h728B, 16'hC556, 16'hCDD7, 16'hC597, 16'hC597, 16'hC597, 16'hB514, 16'hC596, 16'hACD3, 16'hA492,
        16'hACD3, 16'hA493, 16'hA492, 16'hB514, 16'h7B4D, 16'h49C7, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC5D7, 16'h4000, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hBCD3, 16'hE619, 16'hDDD8, 16'hC514, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hB451, 16'hF71C, 16'hFFDF, 16'hFF1E,
        16'hFF1D, 16'hEE9B, 16'hE61A, 16'hD557, 16'hD597, 16'hEE9B, 16'hEE9C, 16'hE65A, 16'hEE5B, 16'hDE1A, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hB452, 16'hCD56, 16'hCD97, 16'hC556, 16'hCD57, 16'hAC52, 16'hA411, 16'hCD57, 16'hCD56, 16'hCD56, 16'hB452, 16'hCD56, 16'hD597, 16'hCD97, 16'hD597, 16'hD597, 16'hCD97, 16'hD598, 16'h9B8E, 16'hC3D1, 16'hED17, 16'hF69C, 16'hFF9F, 16'hEEDC, 16'hA38F, 16'hDDD8, 16'hDD57, 16'h92CD, 16'h928B, 16'hCD16, 16'hDD98, 16'hD597, 16'hD597, 16'hD597, 16'hDD98, 16'hAB8F, 16'hCD15, 16'hD597, 16'hD557, 16'hD557, 16'hD557, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hD598, 16'hD598, 16'hD598, 16'hD5D8, 16'hD598, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hE5D9, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDD97, 16'hA28B, 16'h9148, 16'hDD57, 16'hE619, 16'hE5D9, 16'hE619, 16'hDD98, 16'hA2CC, 16'hED16, 16'hF69C, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFEDD, 16'hF599, 16'hCC94, 16'hAB8F, 16'hEDD8,
        16'hDD97, 16'hEE1A, 16'hE619, 16'hEDD9, 16'hA30D, 16'hE557, 16'hF5D9, 16'hCC12, 16'h930D, 16'hE5D8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hD5D8, 16'hDDD8, 16'hD598, 16'hD598, 16'hDD97, 16'h92CC, 16'hC453, 16'hA38F, 16'hC556, 16'hE65B, 16'hE65A, 16'hE65B, 16'hE65A, 16'hE65B, 16'hE65B, 16'hE65A, 16'hE65B, 16'hE65A, 16'hE65A, 16'hDE19, 16'hDDD9, 16'hDDD9, 16'hD5D8, 16'hD5D9, 16'hD5D8, 16'hDE59, 16'hE69A, 16'hDDD8, 16'h934D, 16'hCD56, 16'hDE19, 16'hDE19, 16'hDE19, 16'h830D, 16'hACD3, 16'hCDD8, 16'hC597, 16'hC597, 16'hC596, 16'hACD3, 16'hBD55, 16'hBD15, 16'hA492, 16'hA493, 16'hA493, 16'hA492, 16'hAD13, 16'h9C51, 16'h000, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9C51, 16'h6A49, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'hBCD3, 16'hEE5B, 16'hD597, 16'hCD56, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD5D7, 16'hCD56, 16'hFFDF, 16'hFF5E, 16'hFF5E, 16'hF6DC, 16'hE65B, 16'hD598, 16'hCD56, 16'hD597, 16'hEE5B, 16'hE65B, 16'hE65A, 16'hEE9B, 16'hDE19, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hCD97, 16'hD597, 16'hD597, 16'hD598, 16'hD598, 16'hB452, 16'hCD56, 16'hCD57, 16'hCD57, 16'hBCD4, 16'hB493, 16'hCD56, 16'hC556, 16'hCD56, 16'hCD56, 16'hAC11, 16'hC556, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'h92CC, 16'hDC94, 16'hED57, 16'hFF1E, 16'hFF9F, 16'hFF5E,
        16'hB412, 16'hDD97, 16'hDD97, 16'hA30E, 16'hAB4E, 16'hBC93, 16'hDDD9, 16'hD598, 16'hD598, 16'hD598, 16'hDDD9, 16'hABD0, 16'hBC52, 16'hDDD8, 16'hD597, 16'hD557, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hE5D9, 16'hE5D9, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hE5D9, 16'hDD97, 16'hA28B, 16'hA20A, 16'hD516, 16'hE61A, 16'hE5D9, 16'hEE1A, 16'hCD15, 16'hAB0E, 16'hF598, 16'hF6DD, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hF61A, 16'hF598, 16'h9ACD, 16'hE557, 16'hDD56, 16'hEE19, 16'hEE1A, 16'hEDD9, 16'hA2CC, 16'hED98, 16'hF6DD, 16'hED98, 16'hA2CC, 16'hBC93, 16'hE619, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'h928B, 16'hCC94, 16'hA38F, 16'hC556, 16'hEE9B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD5D8, 16'hDE19, 16'hE69B, 16'hE619, 16'h9B8E, 16'hC556, 16'hDE19,
        16'hD619, 16'hDE1A, 16'h9BD0, 16'h9C11, 16'hCDD7, 16'hC597, 16'hCDD7, 16'hC597, 16'hACD3, 16'hACD3, 16'hBD55, 16'hA492, 16'hA493, 16'hA492, 16'hA492, 16'hA4D3, 16'hACD2, 16'h4986, 16'h5A89, 16'hF79D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h6A49, 16'hA492, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hC4D4, 16'hEE5A, 16'hC515, 16'hCD97, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hABD0, 16'hF71D, 16'hFFDF, 16'hFF5E, 16'hFF5E, 16'hEE9B, 16'hDE1A, 16'hC515, 16'hCD56, 16'hCD57, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hD5D8, 16'hD598, 16'hD598, 16'hD598, 16'hD597, 16'hD597, 16'hD598, 16'hD598, 16'hD598, 16'hD5D8, 16'hD598, 16'hB453, 16'hCD56, 16'hCD57, 16'hCD56, 16'hC515, 16'hCD56, 16'hC556, 16'hCD56, 16'hCD56, 16'hCD16, 16'hAB8F, 16'hCD56, 16'hD598, 16'hD597, 16'hD597, 16'hD597, 16'hD598, 16'hCD15, 16'hA2CC, 16'hED16, 16'hEDD9, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hBCD4, 16'hC493, 16'hE5D9, 16'hA34E, 16'hC411, 16'hAB4F, 16'hE5D8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'hE619, 16'hBC93, 16'hA30E, 16'hDD98, 16'hD598, 16'hD598, 16'hD598, 16'hD598, 16'hD598, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD8, 16'hDDD9, 16'hE5D9, 16'hE619, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE619, 16'hDD57, 16'hB2CD, 16'hB2CD, 16'hCCD4, 16'hEE5A, 16'hE5D9, 16'hEE1A, 16'hB3D1,
        16'hC3D1, 16'hF619, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFEDD, 16'hFDDA, 16'hC3D1, 16'hC411, 16'hD4D4, 16'hE5D9, 16'hEE1B, 16'hE598, 16'hAB0D, 16'hF5D9, 16'hFF5E, 16'hF6DC, 16'hDCD5, 16'h92CC, 16'hDD98, 16'hE619, 16'hDDD9, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hE5D8, 16'h9ACC, 16'hD4D4, 16'hAB8F, 16'hC556, 16'hEE9C, 16'hE69B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE69B, 16'hE65B, 16'hE69B, 16'hE65B, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD619, 16'hD5D9, 16'hDE19, 16'hE65B, 16'hE65A, 16'h9B8F, 16'hB4D4, 16'hDE1A, 16'hD619, 16'hDE5A, 16'hAC93, 16'h834E, 16'hCDD7, 16'hC597, 16'hC5D7, 16'hC596, 16'hACD3, 16'hA492, 16'hBD15, 16'hA492, 16'hA4D2, 16'hA4D3, 16'hA4D3, 16'hA4D3, 16'hA4D3, 16'h6ACB, 16'h1000, 16'hC5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h3800, 16'hCDD8, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE19, 16'hCD15, 16'hE619, 16'hBCD3, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD5D7, 16'hCD56, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF71D, 16'hE65B, 16'hD597, 16'hC4D5, 16'hCD16, 16'hCD56, 16'hE65A, 16'hE65A, 16'hE65B, 16'hE61A, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD598, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hB453, 16'hCD56, 16'hCD97, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD16, 16'hA34E, 16'hCD56,
        16'hD5D8, 16'hD598, 16'hD597, 16'hD597, 16'hDDD8, 16'hB412, 16'hBBD0, 16'hF598, 16'hF69B, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hDDD9, 16'hA34E, 16'hF61A, 16'hAB4E, 16'hCC94, 16'hA30D, 16'hDD97, 16'hDDD9, 16'hDDD8, 16'hDDD8, 16'hE619, 16'hD516, 16'h9209, 16'hD556, 16'hDDD9, 16'hDDD8, 16'hDD98, 16'hDD98, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hDDD9, 16'hE5D9, 16'hE619, 16'hE61A, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hEE1A, 16'hD4D5, 16'hBB0F, 16'hC390, 16'hC453, 16'hEE5A, 16'hE619, 16'hEE19, 16'hA30D, 16'hDCD5, 16'hF65B, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFEDC, 16'hED58, 16'hAACC, 16'hBB8F, 16'hDD57, 16'hF65B, 16'hDD57, 16'hAB4E, 16'hFE1A, 16'hFF5E, 16'hFF9F, 16'hF619, 16'hB38F, 16'hB412, 16'hEE1A, 16'hDDD9, 16'hDE19, 16'hDDD9, 16'hDDD8, 16'hDDD8, 16'hE5D8, 16'h928C, 16'hD4D5, 16'hAB8F, 16'hC556, 16'hEE9C, 16'hE65B, 16'hE69B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hEE9B,
        16'hE69B, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE65A, 16'hEE5B, 16'hA410, 16'hAC93, 16'hDE5A, 16'hDE19, 16'hDE1A, 16'hCD56, 16'h7B0C, 16'hC597, 16'hC5D7, 16'hC597, 16'hC596, 16'hACD3, 16'hA492, 16'hB4D4, 16'hAC92, 16'hA492, 16'hA4D3, 16'hA4D3, 16'hACD3, 16'hACD3, 16'h838E, 16'h3986, 16'h83CE, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB514, 16'h4801, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDDD8, 16'hCCD5, 16'hDD98, 16'hC4D4, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hABD0, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hEE9B, 16'hE65A, 16'hBC94, 16'hCD16, 16'hB493, 16'hD597, 16'hE69B, 16'hDE5A, 16'hE65A, 16'hD5D8, 16'hD5D8, 16'hDE19, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D9, 16'hD5D9, 16'hD5D8, 16'hB452, 16'hC515, 16'hCD97, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD57, 16'hCD16, 16'h928C, 16'hD557, 16'hD5D8, 16'hD598, 16'hDDD8, 16'hD598, 16'hDDD8, 16'hA34E, 16'hD494, 16'hF598, 16'hFF1D, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hF6DD, 16'hA30D, 16'hEDD9, 16'hB390, 16'hD516, 16'hBC11, 16'hBC52, 16'hE619, 16'hDDD9, 16'hDDD9, 16'hE619, 16'hE5D8, 16'h9209, 16'hBC11, 16'hE619, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD9, 16'hDDD9, 16'hE5D9, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE61A, 16'hE61A, 16'hE5D9, 16'hE5D9, 16'hE5D9,
        16'hE619, 16'hE619, 16'hE619, 16'hEE5A, 16'hC453, 16'hC3D1, 16'hD453, 16'hC452, 16'hEE5A, 16'hE619, 16'hE597, 16'hB2CC, 16'hED98, 16'hF6DC, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFE5B, 16'hD412, 16'hA208, 16'hBC52, 16'hFE5B, 16'hC453, 16'hBBD1, 16'hFE5B, 16'hFF5E, 16'hFF9F, 16'hFEDD, 16'hED57, 16'h928C, 16'hDD97, 16'hE619, 16'hE619, 16'hE619, 16'hDDD8, 16'hDDD8, 16'hDD97, 16'h924B, 16'hD4D5, 16'hABD0, 16'hCD56, 16'hEE9C, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hDE1A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE65A, 16'hEE9B, 16'hB452, 16'hAC52, 16'hE65A, 16'hDE19, 16'hDE1A, 16'hD5D8, 16'h72CB, 16'hBD55, 16'hCDD7, 16'hC597, 16'hBD96, 16'hA4D3, 16'hA492, 16'hAC93, 16'hB4D3, 16'hA451, 16'hACD3, 16'hA4D3, 16'hACD3, 16'hAD14, 16'h9410, 16'h3945, 16'h7BCE, 16'hAD14, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h8B8F, 16'h834E, 16'hFF9F,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD596, 16'hC494, 16'hCCD4, 16'hC556, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC515, 16'hD618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF6DC, 16'hE65A, 16'hD598, 16'hB452, 16'hCD56, 16'hAC11, 16'hDE19, 16'hE65A, 16'hE65A, 16'hE65A, 16'hCD97, 16'hDDD9, 16'hDE19, 16'hDDD9, 16'hD5D8, 16'hD5D8, 16'hDDD9, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD9,
        16'hBC93, 16'hC515, 16'hCD97, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD56, 16'hCD56, 16'hD597, 16'hCD15, 16'h8209, 16'hD597, 16'hDDD8, 16'hD5D8, 16'hDDD8, 16'hDDD8, 16'hDD98, 16'h9B0D, 16'hED56, 16'hEDD9, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hB452, 16'hCC94, 16'hCC53, 16'hCC94, 16'hE597, 16'h9ACC, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hAB4E, 16'hA28B, 16'hE598, 16'hE619, 16'hDDD9, 16'hE5D9, 16'hE5D9, 16'hE5D9, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hE5D9, 16'hE5D9, 16'hE61A, 16'hE619, 16'hE61A, 16'hE61A, 16'hEE5A, 16'hB390, 16'hD494, 16'hDCD5, 16'hBBD0, 16'hEE1A, 16'hEE1A, 16'hD494, 16'hCB90, 16'hF5DA, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF1E, 16'hF5D9, 16'hAA4A, 16'h9B0D, 16'hF5D9, 16'hAB0D, 16'hDCD5, 16'hFE9C, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFE9B, 16'hC412, 16'hA38F, 16'hEE19, 16'hDE19, 16'hDE19, 16'hDDD8, 16'hE619, 16'hDD97, 16'h9209, 16'hDD15,
        16'hB3D0, 16'hCD56, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE65A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE65A, 16'hEE9B, 16'hBCD3, 16'hA411, 16'hDE1A, 16'hDE19, 16'hDE19, 16'hDE19, 16'h7B0C, 16'hACD3, 16'hCDD7, 16'hC597, 16'hC596, 16'hA493, 16'hA492, 16'hA451, 16'hB4D4, 16'h9C51, 16'hACD3, 16'hA4D3, 16'hA4D3, 16'hACD3, 16'hA4D3, 16'h3104, 16'h7BCE, 16'h8C0F, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h6187, 16'hBD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hC514, 16'hBC11, 16'hBC52, 16'hD5D8, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'hB451, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hE65A, 16'hE65A, 16'hB493, 16'hBCD4, 16'hBCD4, 16'hAC11, 16'hE65A, 16'hDE5A, 16'hE65A, 16'hE61A, 16'hCD56, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD5D9, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hC4D4, 16'hC515, 16'hD597, 16'hCD97, 16'hCD57, 16'hCD56, 16'hCD56, 16'hCD57, 16'hD597, 16'hC4D4, 16'h7946, 16'hD557, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hE619, 16'hCD15, 16'hAB0E, 16'hED97, 16'hEE5B, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hE61A, 16'hAB0E, 16'hD494, 16'hC412, 16'hFE5B, 16'hAACD, 16'hD515, 16'hEE5A, 16'hE619, 16'hE619, 16'hEE19, 16'hC452, 16'hA1CA, 16'hC452, 16'hEE1A, 16'hE619, 16'hE619, 16'hE619, 16'hE619,
        16'hE61A, 16'hE619, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hEE5A, 16'hE5D8, 16'hE5D9, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hAB0E, 16'hDD16, 16'hE557, 16'hB34F, 16'hEE1A, 16'hEE5A, 16'hBB8F, 16'hDCD5, 16'hF69B, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF1D, 16'hDCD5, 16'hA30D, 16'hD494, 16'hA2CC, 16'hF5D9, 16'hFF1E, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF1E, 16'hF5D9, 16'h9A4B, 16'hCD15, 16'hE61A, 16'hE5D9, 16'hDDD9, 16'hE619, 16'hDD97, 16'h924A, 16'hDD16, 16'hAB4E, 16'hCD97, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE65A, 16'hEE9B, 16'hBCD4, 16'hA411, 16'hDE5A, 16'hDE19, 16'hDE19, 16'hE65A, 16'h938F, 16'h9C11, 16'hCDD7, 16'hC597, 16'hBD96, 16'hA492, 16'hA492, 16'h9C10, 16'hB493, 16'h9C11, 16'hA4D3, 16'hACD3, 16'hACD3, 16'hACD3, 16'hAD13, 16'h730C, 16'h39C6,
        16'h9CD2, 16'h9450, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD619, 16'h5083, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hBC93, 16'hB3D0, 16'hBC93, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBCD4, 16'hDE19, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hEE5B, 16'hE65A, 16'hDDD8, 16'h9B8F, 16'hCD97, 16'hA3D0, 16'hBC93, 16'hE65A, 16'hDE5A, 16'hE65A, 16'hD5D8,
        16'hCD56, 16'hDE5A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE1A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE61A, 16'hC4D4, 16'hC4D5, 16'hD597, 16'hD597, 16'hCD97, 16'hCD57, 16'hD557, 16'hD597, 16'hDDD8, 16'hBC53, 16'h6800, 16'hD557, 16'hDE19, 16'hDDD9, 16'hDE19, 16'hE61A, 16'hBC52, 16'hC3D1, 16'hED98, 16'hF6DD, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hBC52, 16'hC3D1, 16'hC453, 16'hFE9C, 16'hD494, 16'hAB0D, 16'hEE19, 16'hE619, 16'hE619, 16'hEE5A, 16'hD4D4, 16'hB30D, 16'hA2CC, 16'hE598, 16'hEE1A, 16'hE619, 16'hE619, 16'hE61A, 16'hE61A, 16'hE65A, 16'hEE5A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hE5D8, 16'hE5D9, 16'hE61A, 16'hEE1A, 16'hE61A, 16'hEE5A, 16'hE5D8, 16'hAACD, 16'hE598, 16'hE5D9, 16'hAB4E, 16'hF65A, 16'hE5D8, 16'hBB4E, 16'hEDD8, 16'hFF1E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hF69B, 16'hBB8F, 16'hA2CC, 16'hD494, 16'hFE9C, 16'hFF9F, 16'hFF5F, 16'hFF5F,
        16'hFF5F, 16'hFF5F, 16'hFE9C, 16'hDC94, 16'h9A8C, 16'hE5D9, 16'hE619, 16'hDDD9, 16'hE619, 16'hD556, 16'h9A8C, 16'hE556, 16'hA30D, 16'hD597, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE65A, 16'hEE9B, 16'hC515, 16'hAC11, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE65A, 16'hAC92, 16'h834D, 16'hCDD7, 16'hC5D7, 16'hC596, 16'hA492, 16'hA492, 16'h9C11, 16'hAC52, 16'hAC92, 16'hA492, 16'hB514, 16'hACD3, 16'hACD3, 16'hB514, 16'h8BD0, 16'h6B0C, 16'h8C51, 16'h8C50, 16'hC5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA492, 16'h830C, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hAC11, 16'h9B0E, 16'hC514, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69B, 16'hAC11, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'hE61A, 16'hE65B, 16'hBCD5, 16'hA411, 16'hCDD7, 16'h930E, 16'hD557, 16'hE65A, 16'hDE5A, 16'hE69B, 16'hCD56, 16'hCD57, 16'hE65A, 16'hE65A, 16'hDE59, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE1A, 16'hE61A, 16'hE61A, 16'hE65A, 16'hE65A, 16'hC4D4, 16'hBC93, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hDDD8, 16'hB3D1, 16'h7000, 16'hD556, 16'hE61A, 16'hDDD9, 16'hDE19, 16'hEE1A, 16'hAB8F, 16'hD494, 16'hF5D9, 16'hFF5E, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hE65A, 16'hAA8B, 16'hC412, 16'hF69B, 16'hEDD9, 16'hA24C,
        16'hD4D5, 16'hEE1A, 16'hE619, 16'hEE1A, 16'hDD56, 16'hBB8F, 16'hC411, 16'hBBD0, 16'hF65A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE5B, 16'hDD98, 16'hE5D9, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE5B, 16'hD516, 16'hB34F, 16'hEE1A, 16'hF69B, 16'hBB8F, 16'hFE5B, 16'hCC93, 16'hD453, 16'hF69B, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF1E, 16'hA28A, 16'hBB4F, 16'hF5D9, 16'hFF5E, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFE1A, 16'hAB0E, 16'hBC52, 16'hEE1A, 16'hDDD9, 16'hE61A, 16'hD515, 16'hA30D, 16'hED57, 16'hA30D, 16'hDDD8, 16'hEEDC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE61A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE65A, 16'hE69B, 16'hCD56, 16'hA3D0, 16'hDE19, 16'hDE1A, 16'hDE19, 16'hDE5A, 16'hBD14, 16'h6A8A, 16'hCDD7, 16'hCDD7, 16'hC596,
        16'hA492, 16'h9C92, 16'h9C51, 16'h9C11, 16'hAC92, 16'h9C51, 16'hB514, 16'hACD4, 16'hAD13, 16'hB514, 16'h9411, 16'h9410, 16'h738D, 16'hA513, 16'h8C0F, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h6A09, 16'hBD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h9BCF, 16'h8249, 16'hD5D7, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBC52, 16'hE69B, 16'hFFDF, 16'hFFDF, 16'hFF5E,
        16'hE65A, 16'hE65A, 16'hE65A, 16'h9B8F, 16'hBCD4, 16'hBD14, 16'h8A8C, 16'hDDD8, 16'hE65A, 16'hDE5A, 16'hE65A, 16'hC4D5, 16'hD5D8, 16'hE69A, 16'hE65A, 16'hDE5A, 16'hE61A, 16'hDE19, 16'hE61A, 16'hE65A, 16'hE61A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hC4D5, 16'hB452, 16'hD598, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hE598, 16'hA34E, 16'h8905, 16'hC493, 16'hE61A, 16'hE619, 16'hE61A, 16'hE5D9, 16'hAB0E, 16'hE516, 16'hF65A, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hC493, 16'hA189, 16'hF69C, 16'hFE9C, 16'hDCD5, 16'hAACD, 16'hEE19, 16'hE619, 16'hE619, 16'hE5D8, 16'hB30E, 16'hE517, 16'hA30D, 16'hDD16, 16'hEE5A, 16'hE61A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hE65A, 16'hEE5B, 16'hDD98, 16'hE5D9, 16'hEE1A, 16'hEE1A, 16'hE61A, 16'hF65B, 16'hCC12, 16'hCC52, 16'hF6DC, 16'hF6DC, 16'hBBD1, 16'hEDD8, 16'hC350, 16'hEDD8, 16'hFF1E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F,
        16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hF71D, 16'hC4D4, 16'hF69B, 16'hFF1E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5F, 16'hFEDD, 16'hED17, 16'h9A8C, 16'hE597, 16'hE619, 16'hEE5A, 16'hCD15, 16'hAB4E, 16'hF598, 16'hA30E, 16'hDDD9, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE65A, 16'hE69B, 16'hCD56, 16'hA410, 16'hDE19, 16'hDE1A, 16'hDE19, 16'hDE5A, 16'hCD96, 16'h6208, 16'hC596, 16'hCDD8, 16'hC596, 16'hA492, 16'h9C51, 16'hA451, 16'h93CF, 16'hAC93, 16'h9C10, 16'hB514, 16'hACD3, 16'hAD14, 16'hB514, 16'hA492, 16'h9C11, 16'h9450, 16'h8C51, 16'h9C92, 16'hAD13, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD619, 16'h5905, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'h8B4D, 16'h7A8A, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE19, 16'hB493, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69B, 16'hE61A, 16'hEE9B, 16'hCD57, 16'h930D, 16'hCD56, 16'hB493, 16'h934E, 16'hE619, 16'hE65A, 16'hE65A, 16'hDE19, 16'hBC93, 16'hDE19, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE1A, 16'hE61A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hEE5B, 16'hCD16, 16'hABD1, 16'hDDD8, 16'hD597, 16'hD597, 16'hD598, 16'hD598, 16'hDDD8, 16'hDD57, 16'h9ACC, 16'hAB0D, 16'hAC11, 16'hEE1A, 16'hDE19, 16'hE65A, 16'hD557, 16'hB34F, 16'hED98, 16'hF6DC, 16'hFF9F,
        16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hB2CD, 16'hDDD8, 16'hFF5F, 16'hF61A, 16'hBB4F, 16'hCC12, 16'hEE5A, 16'hE619, 16'hEE5A, 16'hC3D1, 16'hD494, 16'hE557, 16'hA2CB, 16'hEE19, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE5B, 16'hE598, 16'hE5D9, 16'hEE5A, 16'hE61A, 16'hEE1A, 16'hEDD9, 16'hB2CD, 16'hE557, 16'hFF5F, 16'hF69C, 16'hC3D1, 16'hCC12, 16'hDCD4, 16'hF6DD, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFE5B, 16'hCC12, 16'hBC11, 16'hEE1A, 16'hEE5A, 16'hCC94, 16'hBB90, 16'hED98, 16'h9ACD, 16'hE61A, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEEDB, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE65A,
        16'hE69B, 16'hCD57, 16'hAC11, 16'hDE19, 16'hDE1A, 16'hDE19, 16'hDE19, 16'hDDD8, 16'h6A8A, 16'hBD15, 16'hCDD8, 16'hBD56, 16'h9C52, 16'h9410, 16'h9C51, 16'h9410, 16'hAC52, 16'h93D0, 16'hACD3, 16'hB514, 16'hAD14, 16'hAD14, 16'hACD3, 16'h9410, 16'hBD95, 16'h5ACA, 16'hB595, 16'h838E, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAC92, 16'h7B0C, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h728A, 16'h728B, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hA34E, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hE65A, 16'hEE5A, 16'hEE5B, 16'hABD1, 16'hA411, 16'hD5D8, 16'hA411, 16'hA3D0, 16'hE65A, 16'hDE59, 16'hE65A, 16'hD597, 16'hBC93, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE1A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65B, 16'hE65A, 16'hEE9B, 16'hCD56, 16'hA30E, 16'hD598, 16'hDDD8, 16'hD598, 16'hDDD8, 16'hDDD8, 16'hDDD9, 16'hCD16, 16'h9A8C, 16'hD452, 16'h9B4E, 16'hEE1A, 16'hDE19, 16'hEE5A, 16'hCC94, 16'hC3D1, 16'hEDD9, 16'hFF1E, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hF6DC, 16'hD515, 16'hFF5E, 16'hFEDD, 16'hED98, 16'hA9CA, 16'hDD16, 16'hEE5A, 16'hEE5A, 16'hDD16, 16'hBB4F, 16'hFE1A, 16'hCC93, 16'hAB8E, 16'hEE5A, 16'hE61A, 16'hEE1A, 16'hEE1A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE1A, 16'hEE5B, 16'hE598, 16'hE5D8, 16'hEE5A, 16'hE61A, 16'hEE5B, 16'hDD56, 16'hB30E, 16'hF65B, 16'hFF9F, 16'hDD97, 16'hC350,
        16'hDCD5, 16'hF65B, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5F, 16'hFF1D, 16'hF599, 16'hAACD, 16'hDD56, 16'hF61A, 16'hBBD1, 16'hCC52, 16'hED57, 16'h9ACD, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE65A, 16'hE69B, 16'hCD57, 16'hAC11, 16'hDE19, 16'hDE5A, 16'hDE19, 16'hDE19, 16'hE619, 16'h830C, 16'hA452, 16'hCDD8, 16'hBD55, 16'h9C92, 16'h9410, 16'h9C92, 16'h9C11, 16'hA451, 16'h9C11, 16'hA492, 16'hB555, 16'hB514, 16'hAD14, 16'hB514, 16'h8B8F, 16'hC596, 16'h7B8E, 16'h8410, 16'hAD55, 16'h9C91, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h72CB, 16'hAC92, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h6208, 16'h8BCF, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC514, 16'hD5D7, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hE69A, 16'hE65A, 16'hEE9B, 16'hDDD9, 16'h8ACC, 16'hC515, 16'hD598, 16'h82CD, 16'hBCD4, 16'hE65A, 16'hDE59, 16'hE65A, 16'hCD15, 16'hBCD5, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hD597, 16'h9A8C, 16'hD597, 16'hDDD8, 16'hD598, 16'hDDD8, 16'hDDD8, 16'hE619,
        16'hC4D4, 16'h9ACC, 16'hED57, 16'h928B, 16'hDD98, 16'hE61A, 16'hEE1A, 16'hBC11, 16'hD493, 16'hF65A, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF71D, 16'hE61A, 16'hFF1D, 16'hFEDC, 16'hDD16, 16'hB24D, 16'hE557, 16'hEE5A, 16'hEDD9, 16'hBB4F, 16'hED98, 16'hFE1A, 16'hBBD0, 16'hBBD0, 16'hF61A, 16'hEE1A, 16'hE61A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5B, 16'hDD97, 16'hCC53, 16'hEE5A, 16'hE65A, 16'hF65B, 16'hC411, 16'hD4D4, 16'hFF1D, 16'hFF5E, 16'hD4D5, 16'hED98, 16'hF65B, 16'hFF5E, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF1E, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFE9C, 16'hD494, 16'hBBD0, 16'hF5D9, 16'hB30E, 16'hE4D4, 16'hE516, 16'hAB90, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hE61A,
        16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE65A, 16'hE69B, 16'hD597, 16'hAC52, 16'hDE5A, 16'hDE5A, 16'hDE5A, 16'hDE19, 16'hE65A, 16'h938F, 16'h8BCF, 16'hD5D8, 16'hBD55, 16'h9451, 16'h9451, 16'h9451, 16'h9C51, 16'h9BD0, 16'hA452, 16'h9C51, 16'hB514, 16'hB514, 16'hAD14, 16'hB514, 16'h9410, 16'hB514, 16'hAD14, 16'h30C1, 16'hB5D6, 16'h840F, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE5A, 16'h5001, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h5145,
        16'h93CF, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65A, 16'hA38F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'hE65A, 16'hE65A, 16'hEE5B, 16'hB452, 16'h934E, 16'hD5D8, 16'hCD97, 16'h724A, 16'hCD56, 16'hE65A, 16'hDE19, 16'hE61A, 16'hB453, 16'hCD56, 16'hE69B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hDDD9, 16'h8A4B, 16'hCD56, 16'hDDD9, 16'hDDD8, 16'hDDD8, 16'hDDD9, 16'hE619, 16'hBC11, 16'hA30D, 16'hF619, 16'hAB8F, 16'hC494, 16'hEE5B, 16'hEE1A, 16'hB38F, 16'hDCD5, 16'hF69B, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hF65A, 16'hD3D2, 16'hBB0E, 16'hE557, 16'hFE9C, 16'hC412, 16'hD495, 16'hF61A, 16'hF61A, 16'hBC11, 16'hAB0D, 16'hEDD8, 16'hF65B, 16'hEE19, 16'hE597, 16'hF65B, 16'hE65A, 16'hE61A, 16'hE61A,
        16'hEE5B, 16'hE597, 16'hB2CD, 16'hE5D9, 16'hEE5A, 16'hE557, 16'hC34F, 16'hF619, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hF69C, 16'hFF1D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hF69C, 16'hEDD9, 16'hED98, 16'hE598, 16'hE598, 16'hE619, 16'hEE5B, 16'hF6DC, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF1E, 16'hF5D9, 16'hB34F, 16'hE515, 16'hBB4F, 16'hF598, 16'hD494, 16'hB411, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD9, 16'hDE5A, 16'hE69B, 16'hD597, 16'hB493, 16'hDE1A, 16'hDE5A, 16'hDE59, 16'hDE19, 16'hE65A, 16'hAC52, 16'h7B0C, 16'hCD97, 16'hB514, 16'h9450, 16'h9450, 16'h9451, 16'hA492, 16'h938F, 16'hAC52, 16'h93D0, 16'hB514, 16'hB514, 16'hAD14, 16'hB554, 16'h9C51, 16'hA452, 16'hC5D8, 16'h51C7, 16'h7BCF, 16'hAD95, 16'h9410, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD54, 16'h6A4A, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h4945, 16'h9410, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hB3D1, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hE65A, 16'hE65A, 16'hEE5A, 16'hDD98, 16'h820A, 16'hB4D4, 16'hDE19, 16'hCD56, 16'h7A8A, 16'hDDD8, 16'hE61A, 16'hDE19, 16'hDE19, 16'hA3D0, 16'hD5D8, 16'hE69B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE65B,
        16'hEE5B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65A, 16'h928C, 16'hBC93, 16'hDE19, 16'hDDD8, 16'hDDD9, 16'hDDD9, 16'hE619, 16'hA34E, 16'hBB90, 16'hF65A, 16'hD556, 16'h9B0C, 16'hEE1A, 16'hEE1A, 16'hB38F, 16'hE556, 16'hF6DC, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF1D, 16'hED98, 16'hDC94, 16'hBB50, 16'hDCD6, 16'hF5D9, 16'hCC12, 16'hF619, 16'hEDD9, 16'hFE1A, 16'hD4D5, 16'hBB8E, 16'hDCD5, 16'hF61A, 16'hE556, 16'hD4D4, 16'hEE1A, 16'hEE5B, 16'hEE1A, 16'hEE5A, 16'hE598, 16'hA9CA, 16'hE556, 16'hEE1A, 16'hC3D1, 16'hE516, 16'hF71D, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hF71E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hF69B, 16'hED98, 16'hE557, 16'hEDD9, 16'hF69B, 16'hF71D, 16'hFF5E, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFE9C, 16'hE4D5,
        16'hB30E, 16'hCC12, 16'hFE19, 16'hBBD0, 16'hC4D4, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hE61A, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD9, 16'hE65A, 16'hE65B, 16'hD597, 16'hBCD3, 16'hDE19, 16'hDE5A, 16'hDE19, 16'hDE19, 16'hE65A, 16'hB4D4, 16'h6A8A, 16'hC596, 16'hACD3, 16'h8C10, 16'h8C10, 16'h9C51, 16'hA492, 16'h8B8F, 16'hA452, 16'h93CF, 16'hAD14, 16'hAD14, 16'hB514, 16'hB514, 16'hA492, 16'h93CF, 16'hD659, 16'h9410, 16'h4945, 16'hAD95, 16'h8C10, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h7ACB, 16'hACD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71B, 16'h5207, 16'h8BCF, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD55, 16'hCD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9B, 16'hE65B, 16'hE65B, 16'hE619, 16'hAC12, 16'h824A, 16'hD5D7, 16'hDE5A, 16'hB4D4, 16'h7A8B, 16'hE619, 16'hDE19, 16'hE65A, 16'hD598, 16'hA3D0, 16'hE619, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65B, 16'hE65A, 16'hE65A, 16'hEE5B, 16'hE65B, 16'hEE5B, 16'hE65B, 16'hEE9B, 16'hEE5A, 16'h9ACD, 16'hABD0, 16'hE619, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hE5D9, 16'h92CC, 16'hCC52, 16'hF65A, 16'hF69C, 16'h91C8, 16'hD556, 16'hEE5A, 16'hB34F, 16'hED97, 16'hFF1D, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFE9C, 16'hF598, 16'hF61A, 16'hC412, 16'hC390, 16'hC391,
        16'hDD57, 16'hFE5C, 16'hF5D9, 16'hFE5B, 16'hF5D9, 16'hCC93, 16'hCC52, 16'hD493, 16'hD412, 16'hC3D0, 16'hE556, 16'hEE19, 16'hF65B, 16'hEDD9, 16'hCB90, 16'hCC11, 16'hCC12, 16'hD494, 16'hF6DC, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF1D, 16'hEE1A, 16'hE598, 16'hEE5A, 16'hFF1E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF1E, 16'hEEDC, 16'hEE9B, 16'hE65A, 16'hE61A, 16'hE65A, 16'hEE9B, 16'hF71D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hE516, 16'hAACD, 16'hED98, 16'hF5D9, 16'hB34F, 16'hD556, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE619, 16'hE65A, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hDE19, 16'hDDD9, 16'hDE19, 16'hDDD8, 16'hE65A, 16'hEE9B, 16'hD597, 16'hC4D4, 16'hDE1A, 16'hDE5A, 16'hDE19, 16'hDE19, 16'hE65A, 16'hC555, 16'h6A49, 16'hC556, 16'hACD3, 16'h83CF, 16'h8C10, 16'h9C51, 16'hA492, 16'h8BCF, 16'hA411, 16'h9BD0, 16'hACD3,
        16'hB515, 16'hAD14, 16'hB514, 16'hACD3, 16'h838E, 16'hCE18, 16'hB514, 16'h728B, 16'h8C10, 16'hAD95, 16'h8BCF, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'h4904, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71B, 16'h51C7, 16'h83CE, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hAB8F, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hE65B, 16'hEE5B, 16'hE61A, 16'hC515, 16'h934E, 16'h9B4E, 16'hDE19, 16'hDE59, 16'hA411, 16'h8B4E, 16'hE619, 16'hDE19,
        16'hE65A, 16'hC515, 16'hAC52, 16'hE65A, 16'hE65A, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65A, 16'hE65A, 16'hEE5B, 16'hE65B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hA34F, 16'h9B4E, 16'hE619, 16'hDDD9, 16'hDDD9, 16'hDE19, 16'hDD98, 16'h928B, 16'hDCD5, 16'hF65A, 16'hFF5F, 16'hD494, 16'hA2CC, 16'hF619, 16'hBBD0, 16'hED98, 16'hFF1E, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hF69B, 16'hF65A, 16'hFEDC, 16'hE5D8, 16'hC412, 16'hAA4C, 16'hF69C, 16'hFF1D, 16'hF65A, 16'hF61A, 16'hFE5A, 16'hEDD9, 16'hCC12, 16'hC3D1, 16'hDCD5, 16'hC3D1, 16'hC390, 16'hD494, 16'hE516, 16'hDC93, 16'hD493, 16'hCC12, 16'hF69C, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFEDD, 16'hEE1A, 16'hF65B, 16'hFF1D, 16'hFF9F, 16'hFFDF, 16'hFF5F, 16'hF69C, 16'hD557, 16'hB3D1, 16'h92CC, 16'h7146, 16'h6000, 16'h5000, 16'h4800, 16'h4800, 16'h5000,
        16'h6988, 16'h938F, 16'hBCD5, 16'hE61A, 16'hFF1E, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hDDD8, 16'hEE9B, 16'hF65B, 16'hED98, 16'h9ACD, 16'hDDD9, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hDDD8, 16'hEE5A, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hDE19, 16'hDDD8, 16'hDDD8, 16'hD5D8, 16'hE61A, 16'hE69B, 16'hD597, 16'hC515, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE5A, 16'hD5D7, 16'h6A49, 16'hB514, 16'hACD3, 16'h83CE, 16'h8C10, 16'h9C91, 16'hA492, 16'h9410, 16'h93D0, 16'hA411, 16'hA492, 16'hB555, 16'hAD14, 16'hAD14, 16'hB514, 16'h838F, 16'hBD56, 16'hCDD7, 16'h9C10, 16'h9C10, 16'hA554, 16'h9491, 16'hCDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA492, 16'h834D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h628A, 16'h6ACA, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hB390, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hEE9B, 16'hE65B, 16'hE65B, 16'hCD56, 16'hB492, 16'h930D, 16'hAC52, 16'hDE19, 16'hD618, 16'h834E, 16'hA3D0, 16'hE65A, 16'hDE19, 16'hE65A, 16'hBCD4, 16'hBC93, 16'hEE9B, 16'hE65A, 16'hE65B, 16'hE65A, 16'hE65B, 16'hEE5B, 16'hE65A, 16'hE65A, 16'hEE5B, 16'hE65B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hABD0, 16'h8A49, 16'hE5D9, 16'hDE19, 16'hDDD9, 16'hE619, 16'hD557, 16'h9ACC, 16'hED56, 16'hF65B, 16'hFF5F, 16'hFEDD, 16'hB34E, 16'hCC93, 16'hCC52, 16'hEDD8, 16'hFF5E, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F,
        16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hF69C, 16'hF65A, 16'hFF5E, 16'hFF9F, 16'hEE5A, 16'hEE1A, 16'hFFDF, 16'hFF9F, 16'hFF1D, 16'hF69C, 16'hF65B, 16'hFE5B, 16'hEE1A, 16'hF61A, 16'hF65B, 16'hEDD8, 16'hD4D4, 16'hCBD1, 16'hBACD, 16'hE557, 16'hF6DD, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hF6DD, 16'hFF1E, 16'hFF9F, 16'hFF9F, 16'hFF1E, 16'hE5D9, 16'hBBD1, 16'h9209, 16'h7000, 16'h5800, 16'h5800, 16'h5042, 16'h50C3, 16'h48C4, 16'h4904, 16'h48C4, 16'h4082, 16'h3000, 16'h2000, 16'h000, 16'h3000, 16'h7A8B, 16'hCD57, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFE9C, 16'hE556, 16'h9ACD, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hDDD8, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hDE19, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hE619, 16'hE69B, 16'hD597, 16'hC515, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19,
        16'hDE18, 16'h7A8B, 16'hACD3, 16'hACD2, 16'h7BCE, 16'h8C50, 16'h9C91, 16'hA492, 16'h9C51, 16'h8B8E, 16'hA452, 16'h9C51, 16'hB554, 16'hAD14, 16'hAD14, 16'hB555, 16'h8C10, 16'hAD14, 16'hD619, 16'hA451, 16'hB4D4, 16'h8C0F, 16'hB595, 16'h940F, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h6208, 16'hC597, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5C, 16'h734C, 16'h4985, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hBC52, 16'hDDD8, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'hE65B,
        16'hE69B, 16'hCD97, 16'hAC92, 16'hBCD4, 16'h82CC, 16'hC515, 16'hDE59, 16'hCD97, 16'h61C8, 16'hAC93, 16'hE61A, 16'hDE19, 16'hE65A, 16'hA3D0, 16'hC515, 16'hEE9B, 16'hE65A, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hEE9B, 16'hC494, 16'h7000, 16'hDD97, 16'hE61A, 16'hDE19, 16'hE61A, 16'hD515, 16'hAB4E, 16'hED97, 16'hF69C, 16'hFF5F, 16'hFF5F, 16'hF65B, 16'hBB0E, 16'hBB4F, 16'hF619, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF1E, 16'hF69C, 16'hF6DD, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hF6DD, 16'hFEDD, 16'hFF1E, 16'hFF5E, 16'hFF1E, 16'hFF1D, 16'hFEDC, 16'hF619, 16'hEDD9, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF5F, 16'hF65C, 16'hCC13,
        16'h90C6, 16'h7000, 16'h7105, 16'h7987, 16'h7187, 16'h6105, 16'h58C4, 16'h58C4, 16'h5083, 16'h4883, 16'h4082, 16'h4082, 16'h4083, 16'h40C4, 16'h4104, 16'h38C4, 16'h000, 16'h2000, 16'h938F, 16'hC515, 16'hEE1A, 16'hDD57, 16'hDD98, 16'hFF9F, 16'hFF9F, 16'hFEDD, 16'hCC53, 16'hA38F, 16'hF69C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hDDD8, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hD598, 16'hDE19, 16'hEE9B, 16'hD597, 16'hCD56, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'h830D, 16'hA492, 16'h9C91, 16'h7BCE, 16'h8C10, 16'h9C51, 16'h9C51, 16'hA452, 16'h834E, 16'hA451, 16'h940F, 16'hB555, 16'hAD14, 16'hAD14, 16'hB555, 16'h9451, 16'h9C92, 16'hD619, 16'hB514, 16'hB514, 16'hBCD4, 16'h9CD2, 16'h9C91, 16'hC5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC5D7, 16'h5187, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h8C0F, 16'h000, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC493, 16'hBC93, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hE69B, 16'hEE9B, 16'hDDD9, 16'hAC93, 16'hB4D4, 16'hC515, 16'h82CC, 16'hD597, 16'hDE19, 16'hBD15, 16'h4883, 16'hB4D4, 16'hE61A, 16'hDE19, 16'hDE19, 16'h9B4E, 16'hD597, 16'hE69B, 16'hE65B, 16'hE65B, 16'hE69B, 16'hE65B, 16'hEE9B, 16'hE65B, 16'hE65A, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hE69B, 16'hEE9C, 16'hD556, 16'h6800, 16'hCCD4, 16'hEE5A, 16'hE619, 16'hEE5A, 16'hC4D4, 16'hB38F, 16'hED98, 16'hF6DD, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hEDD9, 16'hA1CA,
        16'hEDD9, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF5F, 16'hFF1D, 16'hF6DD, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hF61B, 16'hDBD2, 16'hA188, 16'h8187, 16'h8187, 16'h8187, 16'h7146, 16'h6146, 16'h5905, 16'h5104, 16'h50C4, 16'h48C4, 16'h48C3, 16'h4904, 16'h4904, 16'h4904, 16'h40C3, 16'h4042, 16'h4042, 16'h40C3, 16'h40C3, 16'h1000, 16'h2800, 16'h6002, 16'hAB0E, 16'hF69C, 16'hFF9F, 16'hFF9F, 16'hFF1D, 16'hB390, 16'hC4D4, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE61A, 16'hDDD8, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hE61A, 16'hD5D8,
        16'hDDD8, 16'hDDD8, 16'hD598, 16'hDE19, 16'hE69B, 16'hD597, 16'hCD56, 16'hDE19, 16'hDE19, 16'hDE5A, 16'hDE5A, 16'hDE19, 16'hDE1A, 16'h938E, 16'h93CF, 16'h9410, 16'h7BCE, 16'h8C10, 16'h9C51, 16'h9C51, 16'hA492, 16'h834E, 16'h9C11, 16'h93CF, 16'hB514, 16'hAD14, 16'hB514, 16'hB514, 16'hA492, 16'h9410, 16'hCE18, 16'hCDD7, 16'hA492, 16'hE65A, 16'h8BD0, 16'hAD95, 16'h8C0F, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h8B8E, 16'hA452, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD14, 16'h000, 16'hAD13, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD597, 16'hB3D0, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'hEE9B, 16'hE65A, 16'hBCD4, 16'hAC93, 16'hC556, 16'hC515, 16'h8B0D, 16'hD5D8, 16'hD5D8, 16'hAC52, 16'h4000, 16'hBD15, 16'hDE19, 16'hDE19, 16'hD5D8, 16'h930D, 16'hDE19, 16'hE69B, 16'hE65B, 16'hE65B, 16'hE69B, 16'hE65B, 16'hEE5B, 16'hE65B, 16'hE65A, 16'hE65B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hE5D9, 16'h7843, 16'hABD0, 16'hEE5A, 16'hDE19, 16'hEE5A, 16'hBC52, 16'hBBD1, 16'hF5D9, 16'hFF1D, 16'hFF5F, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hEDD9, 16'hE619, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF1E, 16'hF69C, 16'hF65B, 16'hEDD9, 16'hF5D9, 16'hEDD9, 16'hF61A, 16'hF69C, 16'hFF1E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFE9D, 16'hDC14, 16'hB20A, 16'h99C8, 16'h89C7, 16'h7987, 16'h6145, 16'h4000, 16'h2000, 16'h1800, 16'h2800, 16'h3800, 16'h3800, 16'h4000, 16'h2000, 16'h000, 16'h000, 16'h2000, 16'h4082, 16'h4904, 16'h48C3, 16'h4882, 16'h50C4, 16'h5945, 16'h48C2, 16'h5104, 16'h82CC, 16'hCD16, 16'hFF1D, 16'hFF1D, 16'h9ACD, 16'hD597, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE5D9, 16'hDDD8, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hDE19, 16'hD5D8, 16'hDDD8, 16'hDDD8, 16'hD598, 16'hDE19, 16'hEE9B, 16'hD5D8, 16'hCD56, 16'hDE19, 16'hDE5A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE65A, 16'hA411, 16'h72CB, 16'h8C10, 16'h840F, 16'h8C0F, 16'h9C51, 16'h9C51, 16'hA492, 16'h8B8F, 16'h9C10, 16'h93CF, 16'hACD3, 16'hB514, 16'hAD14, 16'hB514, 16'hA4D3, 16'h8C0F, 16'hC5D7, 16'hD618, 16'h9C50, 16'hE69A, 16'hC556, 16'h9491, 16'h9491, 16'hC5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'h50C5, 16'hDE5A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE58, 16'h1000, 16'h83CE, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE19, 16'hAB4E, 16'hFF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hEE9B, 16'hE65A, 16'hC515, 16'hAC93, 16'hB4D3, 16'hDE18, 16'hCD56, 16'h938F, 16'hD5D8, 16'hCD56, 16'h9BCF, 16'h5146, 16'hC556, 16'hDE19, 16'hDE5A, 16'hCD56, 16'h934E, 16'hE65A, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hE61A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hEE5A, 16'h8A09, 16'h8A4A,
        16'hE619, 16'hE619, 16'hEE5A, 16'hB411, 16'hCC53, 16'hF5D9, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF1D, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hF6DC, 16'hF65B, 16'hF65A, 16'hEE1A, 16'hEE1A, 16'hEDD9, 16'hEDD9, 16'hED97, 16'hE557, 16'hF5D9, 16'hFEDC, 16'hFF5E, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF1D, 16'hDCD6, 16'hC2CE, 16'hAA4B, 16'h89C8, 16'h78C4, 16'h5800, 16'h5000, 16'h7A09, 16'hAC52, 16'hCD56, 16'hD5D8, 16'hDE19, 16'hE65A, 16'hE65A, 16'hDDD9, 16'hCD97, 16'hB4D3, 16'h830D, 16'h4000, 16'h000, 16'h3800, 16'h5105, 16'h5083, 16'h4000, 16'h5105, 16'h5905, 16'h4000, 16'h4800, 16'hBC12, 16'hED98, 16'h928B, 16'hEE5A, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B,
        16'hEE9B, 16'hDDD8, 16'hE619, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hDDD9, 16'hD5D8, 16'hD598, 16'hD598, 16'hD597, 16'hE61A, 16'hEE9B, 16'hD5D8, 16'hCD56, 16'hDE19, 16'hDE19, 16'hE61A, 16'hDE19, 16'hDE19, 16'hE65A, 16'hAC52, 16'h6ACA, 16'h8C10, 16'h840F, 16'h8C0F, 16'h9C91, 16'h9C51, 16'h9C92, 16'h8BCF, 16'h93CF, 16'h938F, 16'hACD3, 16'hB514, 16'hAD14, 16'hB514, 16'hAD13, 16'h838E, 16'hC596, 16'hD619, 16'hB514, 16'hB555, 16'hF75D, 16'h8BCF, 16'hAD54, 16'h8C10, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'h9411, 16'h8B8F, 16'hFFDE, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h5A8A, 16'h5A49, 16'hDE9A, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'h9ACC, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'hEE5B, 16'hC516, 16'hAC52, 16'hAC93, 16'hC556, 16'hE65A, 16'hC515, 16'h9BD0, 16'hD5D8, 16'hAC92, 16'h8B8F, 16'h59C7, 16'hCD56, 16'hDE19, 16'hE65A, 16'hBCD4, 16'h9B8F, 16'hE65B, 16'hE65A, 16'hE65B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE61A, 16'hE65B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hA34E, 16'h7000, 16'hDD97, 16'hE65A, 16'hEE5A, 16'hB38F, 16'hD494, 16'hF61A, 16'hFF5E, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF1D, 16'hF69C, 16'hF6DC, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hF69C, 16'hDC13, 16'hB28C, 16'hA20A, 16'hA0C7, 16'h91C9, 16'hBC93, 16'hE61A, 16'hFF1D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF5F, 16'hFF5E, 16'hFF1E, 16'hE65B, 16'hBCD4, 16'h724A, 16'h2800, 16'h5843, 16'h71C8, 16'h4000, 16'h3000, 16'h5802, 16'h6987, 16'h8209, 16'h9189, 16'hBC11, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hDD97, 16'hE619, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hDDD8, 16'hD5D8, 16'hE65A, 16'hEE9B, 16'hDDD8, 16'hCD56, 16'hDDD9, 16'hDE19, 16'hDE1A, 16'hDE1A, 16'hDE19, 16'hE65A, 16'hB493, 16'h72CA, 16'h8C0F, 16'h840F, 16'h8C0F, 16'h9C91, 16'h9C92, 16'h9C92, 16'h9410, 16'h8B8F, 16'h9BCF, 16'hA492, 16'hB555, 16'hB514, 16'hB514, 16'hB514, 16'h7B8E, 16'hBD55, 16'hCE18,
        16'hCDD8, 16'h9410, 16'hFF9E, 16'hC596, 16'h9C91, 16'h9491, 16'hC5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h5186, 16'hCDD8, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDE, 16'h9450, 16'h3103, 16'hBD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'h9B4D, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5D, 16'hEE9B, 16'hD597, 16'hAC52, 16'hAC52, 16'hC515, 16'hDE19, 16'hE65A, 16'hCD16, 16'hA3D0, 16'hD597, 16'h9C10, 16'h8BCF, 16'h59C8, 16'hCD97, 16'hDE19, 16'hE65A, 16'hAC52, 16'hAC52, 16'hEE9B, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B,
        16'hEE5B, 16'hEE9B, 16'hE619, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hBC53, 16'h8000, 16'hBC52, 16'hEE5A, 16'hEE5A, 16'hB38F, 16'hDCD5, 16'hF65B, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF1E, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hF69C, 16'hDC54, 16'hCB91, 16'hD3D2, 16'hD516, 16'hF71D, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hFF5E, 16'hFF5F, 16'hFEDD, 16'hCD16, 16'h7105, 16'hCC93,
        16'hE5D9, 16'hB412, 16'h8A8B, 16'h68C4, 16'hA2CC, 16'h9188, 16'hCD15, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE9C, 16'hE61A, 16'hD557, 16'hEE5A, 16'hEEDC, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE5B, 16'hD5D8, 16'hDDD8, 16'hD598, 16'hE61A, 16'hDDD9, 16'hE65A, 16'hEE9B, 16'hDDD8, 16'hCD56, 16'hD5D8, 16'hDE19, 16'hDE1A, 16'hDE5A, 16'hDE19, 16'hE65A, 16'hBD14, 16'h6A49, 16'h8C0F, 16'h8C0F, 16'h8C0F, 16'h9451, 16'h9C51, 16'h9C51, 16'h9451, 16'h8B8E, 16'h9BD0, 16'h9C51, 16'hB555, 16'hAD14, 16'hB514, 16'hB515, 16'h7B8E, 16'hACD3, 16'hCE18, 16'hD618, 16'h9C51, 16'hD659, 16'hFF9E, 16'h8BCE, 16'hA554, 16'h8BCF, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD14, 16'h72CC, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE18, 16'h4A07, 16'h8C0F, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'h9B4D, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hEE9B, 16'hDE19, 16'hB493, 16'hAC52, 16'hB4D4, 16'hD5D8, 16'hDE19, 16'hDE19, 16'hCD56, 16'hA3D0, 16'hB4D3, 16'h8BCF, 16'h9410, 16'h6208, 16'hCD96, 16'hDE19, 16'hE65A, 16'h938F, 16'hC4D4, 16'hEE9B, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE61A, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF69C, 16'hCD16, 16'h8946, 16'h9ACC, 16'hE5D9, 16'hEE5A, 16'hB38E, 16'hE516, 16'hF65B, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hF71D, 16'hDE19, 16'hC4D4, 16'hAB90, 16'h92CD, 16'h92CC, 16'h924B, 16'h924B, 16'hAB0E, 16'hCC12, 16'hED57, 16'hF65B, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF5E, 16'hF65C, 16'hEE1A, 16'hF6DD, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFEDD, 16'hFEDD, 16'hFF1D, 16'hFF1E, 16'hFF1E, 16'hEE5A, 16'hB3D1, 16'hEDD9, 16'hFF1E, 16'hFEDC, 16'hE61A, 16'hCCD5, 16'hAACC, 16'hEE1A, 16'hF69C, 16'hEE9B, 16'hE65A, 16'hEE5B, 16'hEE9C, 16'hE5D9, 16'hD597, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hE65A, 16'hD598, 16'hDDD9, 16'hD598, 16'hE61A, 16'hDDD9, 16'hE65A, 16'hEE9B, 16'hDDD8, 16'hCD16, 16'hCD97, 16'hDE19, 16'hDE5A, 16'hDE5A, 16'hDE5A, 16'hE65A, 16'hC515, 16'h6248, 16'h8C0F, 16'h8C0F, 16'h8C0F, 16'h9451, 16'h9C51,
        16'h9C51, 16'h9C51, 16'h8B8E, 16'h9C10, 16'h93D0, 16'hB554, 16'hAD14, 16'hAD14, 16'hB555, 16'h83CF, 16'hA492, 16'hCDD8, 16'hCE18, 16'hBD55, 16'hAD13, 16'hFFDF, 16'hBD56, 16'h9CD1, 16'h8C50, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h6208, 16'hCDD8, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h734D, 16'h5289, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'h9B0D, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hDE59, 16'hDE19, 16'hC516, 16'hAC52, 16'hAC93, 16'hCD97, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD598, 16'h9B8F, 16'h9BD0, 16'h9410, 16'h8BCF,
        16'h6208, 16'hCD96, 16'hDE5A, 16'hDE19, 16'h7A8B, 16'hCD56, 16'hEE9B, 16'hE65B, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE61A, 16'hE61A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hDDD8, 16'h9A4A, 16'h9A09, 16'hD556, 16'hEE5A, 16'hAB4E, 16'hE556, 16'hF65B, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hEE9B, 16'hB493, 16'h7A09, 16'h5000, 16'h4800, 16'h5000, 16'h5800, 16'h6003, 16'h7105, 16'h8187, 16'h89C8, 16'h9188, 16'hA20A, 16'hC38F, 16'hDD15, 16'hF6DD, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1D, 16'hFF1D,
        16'hFF1D, 16'hFEDD, 16'hFEDD, 16'hFEDD, 16'hFEDD, 16'hFEDD, 16'hFEDC, 16'hFEDD, 16'hFEDD, 16'hFEDC, 16'hFF1D, 16'hF65B, 16'hE598, 16'hF65B, 16'hF69B, 16'hFEDD, 16'hEDD9, 16'hA38F, 16'hF6DC, 16'hEEDC, 16'hEE5B, 16'hE619, 16'hEE9B, 16'hEE9C, 16'hDDD8, 16'hDD97, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hDE19, 16'hDDD8, 16'hE65A, 16'hD598, 16'hDDD9, 16'hD5D8, 16'hE65A, 16'hEE9B, 16'hDDD9, 16'hCD16, 16'hCD56, 16'hDE19, 16'hE65A, 16'hDE5A, 16'hDE19, 16'hE65A, 16'hC515, 16'h6249, 16'h8C10, 16'h8C0F, 16'h8C0F, 16'h9451, 16'h9C51, 16'h9C51, 16'h9C92, 16'h8B8E, 16'hA410, 16'h93D0, 16'hB555, 16'hAD14, 16'hAD14, 16'hB555, 16'h9410, 16'h9451, 16'hCDD7, 16'hCDD8, 16'hC5D7, 16'h8BCF, 16'hF79E, 16'hEF1C, 16'h83CF, 16'hA513, 16'hA4D2, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB514, 16'h7ACC, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB595, 16'h4A48, 16'h8C0F, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'hA34E, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hCD55, 16'hBC93, 16'hD5D8, 16'hAC93, 16'hA452, 16'hC555, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD9, 16'h9BD0, 16'h8BCF, 16'h9411, 16'h93D0, 16'h6208, 16'hC556, 16'hDE19, 16'hD5D8, 16'h724A, 16'hDDD9, 16'hEE9B, 16'hE65B, 16'hE69B, 16'hE65B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hDDD9, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE1A, 16'h9ACC, 16'hAA8D, 16'hB412, 16'hF65A, 16'hAB0D, 16'hE557, 16'hF69C, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF1E, 16'hC515, 16'h5842, 16'h3800, 16'h4800, 16'h5905, 16'h6146, 16'h6947,
        16'h6946, 16'h7146, 16'h7987, 16'h81C8, 16'h89C8, 16'h9209, 16'h9A09, 16'hAA0A, 16'hBACD, 16'hCC12, 16'hEE5B, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFEDD, 16'hFEDD, 16'hFEDD, 16'hFEDD, 16'hFEDD, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFEDC, 16'hFE9C, 16'hF65B, 16'hFE5B, 16'hBC11, 16'hCCD4, 16'hFF1D, 16'hEE9C, 16'hE61A, 16'hE619, 16'hEE9C, 16'hEE9B, 16'hDD57, 16'hDDD8, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEE9C, 16'hDDD8, 16'hDE19, 16'hEE5B, 16'hDDD8, 16'hD598, 16'hD597, 16'hE65A, 16'hEE9B, 16'hDE19, 16'hCD16, 16'hBCD5,
        16'hD5D8, 16'hE65A, 16'hDE19, 16'hDE19, 16'hE65A, 16'hC515, 16'h6248, 16'h8C0F, 16'h8C0F, 16'h8C0F, 16'h9451, 16'h9C51, 16'h9C51, 16'hA492, 16'h838E, 16'hA410, 16'h8B8F, 16'hB554, 16'hAD14, 16'hAD14, 16'hB555, 16'h9C51, 16'h83CF, 16'hC5D7, 16'hC5D7, 16'hCE18, 16'h9410, 16'hD69A, 16'hFFDF, 16'hA492, 16'h9D13, 16'h840F, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DC, 16'h5945, 16'hD618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C0F, 16'h6B8D, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE699, 16'hB411, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5D, 16'hBC52, 16'h9B4E, 16'hCD57, 16'hBCD4,
        16'h9C10, 16'hB4D4, 16'hD619, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD619, 16'hDE19, 16'hA3D0, 16'h7B0C, 16'h9C51, 16'h8BCF, 16'h59C7, 16'hC556, 16'hE65A, 16'hCD56, 16'h7A8A, 16'hE65A, 16'hEE9B, 16'hE65B, 16'hE69B, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hDDD8, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hA38E, 16'hC350, 16'h9A8C, 16'hE598, 16'hBB90, 16'hE557, 16'hF6DD, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1D, 16'hA3D0, 16'h3000, 16'h4883, 16'h5105, 16'h50C4, 16'h58C4, 16'h6105, 16'h6105, 16'h6146, 16'h6145, 16'h60C3, 16'h6001, 16'h6800, 16'h7002, 16'h88C5, 16'hA209, 16'hBACD, 16'hD391, 16'hE4D5, 16'hF6DC, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F,
        16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF6DC, 16'hFEDD, 16'hFE9C, 16'hFE9C, 16'hFEDD, 16'hFE9C, 16'hF65B, 16'hFE9C, 16'hF65B, 16'hF69C, 16'hFE9C, 16'hF69C, 16'hF65B, 16'hF65B, 16'hF69C, 16'hFE9C, 16'hF65B, 16'hF65B, 16'hF61B, 16'hA2CD, 16'hE619, 16'hF6DC, 16'hF69C, 16'hDDD8, 16'hEE5B, 16'hF69C, 16'hEE5A, 16'hD516, 16'hE5D9, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hEE5B, 16'hDD98, 16'hE61A, 16'hEE5B, 16'hD598, 16'hD598, 16'hD598, 16'hE65A, 16'hE69B, 16'hDE19, 16'hCD15, 16'hBCD4, 16'hD5D8, 16'hE65A, 16'hDE1A, 16'hDE19, 16'hDE1A, 16'hCD56, 16'h6A49, 16'h940F, 16'h8C10, 16'h8C0F, 16'h9450, 16'h9451, 16'h9C51, 16'hA492, 16'h838E, 16'h9C10, 16'h8B8E, 16'hB554, 16'hAD14, 16'hAD14, 16'hB554, 16'hA492, 16'h838E, 16'hC5D7, 16'hC5D8, 16'hCE19, 16'hA4D3, 16'hB555, 16'hFFDF, 16'hDE5A, 16'h8C50, 16'h94D2, 16'hB555, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9C52,
        16'h8B8E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE18, 16'h6B4C, 16'h844F, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'hA30D, 16'hF6DC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hB411, 16'hABD0, 16'hBD15, 16'hD597, 16'hA411, 16'hA452, 16'hCD97, 16'hDE5A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD5D8, 16'hD618, 16'hBCD4, 16'h6A8A, 16'h9410, 16'h8BCF, 16'h6208, 16'hCD56, 16'hE65A, 16'hBCD4, 16'h830C, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hDD98, 16'hEE5A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF69C, 16'hBC52, 16'hBB0F, 16'hC3D1, 16'hB38F, 16'hC3D1, 16'hE556, 16'hFF1D, 16'hFF9F, 16'hFF5E,
        16'hFF5E, 16'hFF9F, 16'hF6DC, 16'h8B0D, 16'h4800, 16'h6146, 16'h4882, 16'h4842, 16'h5083, 16'h5905, 16'h5104, 16'h3800, 16'h3800, 16'h4800, 16'h6000, 16'h7986, 16'h8A0A, 16'h924A, 16'h9A0A, 16'hAA4B, 16'hBACC, 16'hCB91, 16'hDCD5, 16'hF6DC, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1E, 16'hFF1D, 16'hFEDD, 16'hFF1D, 16'hFEDC, 16'hFEDD, 16'hFEDD, 16'hF69C, 16'hFE9C, 16'hFE9C, 16'hF65B, 16'hFE9C, 16'hF65B, 16'hF65B, 16'hF69C, 16'hFE9C, 16'hF65A, 16'hF61B, 16'hFE5C, 16'hFE9C, 16'hF61A, 16'hF65B, 16'hFE5B, 16'hDD15, 16'hA30E, 16'hFEDC, 16'hF6DC, 16'hE61A, 16'hD597, 16'hF69C, 16'hF69C, 16'hE619, 16'hD556, 16'hE61A, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEEDC,
        16'hE65A, 16'hDDD8, 16'hE61A, 16'hE65B, 16'hD598, 16'hDD98, 16'hDDD8, 16'hE65A, 16'hEE9B, 16'hE619, 16'hC515, 16'hB493, 16'hCD97, 16'hE65A, 16'hDE1A, 16'hDE19, 16'hDE1A, 16'hCD57, 16'h6A49, 16'h9410, 16'h8C50, 16'h8C0F, 16'h9410, 16'h9451, 16'h9C91, 16'hA493, 16'h838F, 16'h9C10, 16'h8B8E, 16'hAD14, 16'hAD14, 16'hAD14, 16'hAD14, 16'hACD3, 16'h7B8E, 16'hBD96, 16'hCDD8, 16'hCE18, 16'hBD97, 16'h9C91, 16'hFFDF, 16'hFF9F, 16'h9C51, 16'h9D53, 16'h840F, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE5A, 16'h50C2, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9C92, 16'h6B8C, 16'h9CD2, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE659, 16'hAB8F,
        16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hABD0, 16'hC515, 16'hC555, 16'hD596, 16'hBCD4, 16'h9C11, 16'hC556, 16'hDE19, 16'hDE5A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hCD97, 16'hD5D8, 16'hCD56, 16'h724A, 16'h8BCF, 16'h93D0, 16'h59C7, 16'hBD15, 16'hE65A, 16'hAC52, 16'h938F, 16'hEE9B, 16'hE65B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hD557, 16'hE61A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF69C, 16'hD556, 16'h9A0B, 16'hED16, 16'hAB4F, 16'hAACD, 16'hED98, 16'hFF1D, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hF6DC, 16'h7A4A, 16'h1800, 16'h5145, 16'h4841, 16'h4001, 16'h50C3, 16'h5104, 16'h3000, 16'h4800, 16'h930C, 16'hBCD4, 16'hDDD8, 16'hEE9B, 16'hF6DC, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF6DC, 16'hF69B, 16'hF65B, 16'hF69C, 16'hFF1E, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFEDD, 16'hFEDD, 16'hFEDD, 16'hFE9C, 16'hFEDD, 16'hF65C, 16'hFE9C, 16'hFE9C, 16'hF65B, 16'hF65C, 16'hF65C, 16'hF5DA, 16'hF61A, 16'hFE9C, 16'hF61A, 16'hF61A, 16'hFE5B, 16'hFE9C, 16'hF5DA, 16'hF65B, 16'hF61B, 16'hFE1B, 16'hBBD1, 16'hCCD5, 16'hFF1D, 16'hF6DC, 16'hD556, 16'hE619, 16'hF69C, 16'hEE9C, 16'hE5D9, 16'hD557, 16'hEE5A, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hE619, 16'hDDD8, 16'hE65A, 16'hE65A, 16'hDDD8, 16'hDDD8, 16'hD5D8, 16'hE65A, 16'hEE9B, 16'hDE19, 16'hC4D5, 16'hB452, 16'hCD56, 16'hE65A, 16'hDE1A, 16'hDE1A, 16'hE61A, 16'hD597, 16'h728A, 16'h8C0F, 16'h8C50, 16'h8C0F, 16'h9450, 16'h9C51, 16'h9C92, 16'hA4D3, 16'h8B8F, 16'h9C10, 16'h8B8E, 16'hAD14, 16'hAD14, 16'hAD14, 16'hB554, 16'hAD14, 16'h734D, 16'hB555, 16'hCE18, 16'hC5D7, 16'hCE18, 16'h8C10, 16'hDE9A, 16'hFFDF, 16'hCDD7, 16'h8C91,
        16'h8490, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h7B0C, 16'hACD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h8C50, 16'h744F, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD618, 16'h9B0C, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'hA34E, 16'hD597, 16'hDE59, 16'hC556, 16'hCD96, 16'h9BD0, 16'hB4D4, 16'hDE19, 16'hDE5A, 16'hDE19, 16'hDE19, 16'hDE5A, 16'hC596, 16'hC556, 16'hD5D8, 16'hD5D9, 16'h938E, 16'h6ACB, 16'h9C11, 16'h5986, 16'hB4D4, 16'hE65A, 16'h938F, 16'hA410, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hE65B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hDD98, 16'hDDD8, 16'hEE9B, 16'hEE9B, 16'hEE9B,
        16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hE619, 16'hA28B, 16'hDCD5, 16'hE557, 16'h920A, 16'hD4D5, 16'hFF5E, 16'hFF5E, 16'hEE9B, 16'hDDD8, 16'h82CC, 16'h3800, 16'h5105, 16'h3800, 16'h4042, 16'h5945, 16'h4000, 16'h4800, 16'hAC11, 16'hE65A, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1E, 16'hFEDD, 16'hFEDD, 16'hFEDD, 16'hFE9C, 16'hFF1D, 16'hFE9C, 16'hFE9C, 16'hFEDC, 16'hF65C, 16'hF65B, 16'hFE9C, 16'hF5DA, 16'hF5D9, 16'hFE9C, 16'hF61B, 16'hF5D9, 16'hF65B, 16'hFE9C, 16'hF5D9, 16'hF65B, 16'hF61B, 16'hF61A, 16'hF5DA, 16'h9ACC, 16'hEE5A, 16'hF6DC, 16'hE61A, 16'hCCD4,
        16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hDDD8, 16'hDD97, 16'hEE5B, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hE619, 16'hE619, 16'hE61A, 16'hE619, 16'hDDD9, 16'hDDD8, 16'hD5D8, 16'hE69B, 16'hEE9B, 16'hDE19, 16'hC4D4, 16'hAC11, 16'hC556, 16'hE65A, 16'hDE1A, 16'hDE1A, 16'hE65A, 16'hCD57, 16'h6208, 16'h9410, 16'h8C10, 16'h8C0F, 16'h9450, 16'h9C91, 16'hA4D2, 16'hACD3, 16'h8BCF, 16'h9C10, 16'h8B8E, 16'hAD14, 16'hAD14, 16'hAD14, 16'hAD14, 16'hAD14, 16'h83CE, 16'hAD14, 16'hCE18, 16'hC5D7, 16'hCE19, 16'hA4D3, 16'hBD96, 16'hFFDF, 16'hF75D, 16'h8C50, 16'h9512, 16'h9C92, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD96, 16'h59C6, 16'hF75C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C50, 16'h7C90, 16'hCE18, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE19, 16'h928B, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'h8A09, 16'hD618, 16'hFF5D, 16'hC515, 16'hDDD8, 16'hB493, 16'hA411, 16'hCD97, 16'hE65A, 16'hDE5A, 16'hDE19, 16'hDE5A, 16'hD5D8, 16'hACD3, 16'hCD97, 16'hD5D8, 16'hD618, 16'hBD14, 16'h5146, 16'h93D0, 16'h6249, 16'hA452, 16'hE619, 16'h82CC, 16'hB493, 16'hEE9B, 16'hE65B, 16'hEE9B, 16'hE65A, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hDDD8, 16'hD557, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hAB4E, 16'hCC13, 16'hEDD9, 16'hEDD8, 16'hDD16, 16'hE5D9, 16'hDD98, 16'hD515, 16'h7946, 16'h3000, 16'h4904, 16'h3000, 16'h40C3, 16'h48C3, 16'h3800, 16'h930D, 16'hE619, 16'hFF5F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1E, 16'hFF1D, 16'hFEDD, 16'hFF1D, 16'hFE9C, 16'hFEDD, 16'hFEDC, 16'hF65B, 16'hFEDD, 16'hFE9C, 16'hF61B, 16'hFE9C, 16'hFE5B, 16'hF5D9, 16'hF65C, 16'hFE5C, 16'hF5D9, 16'hF61A, 16'hFE5C, 16'hF5D9, 16'hFE5B, 16'hF5DA, 16'hF5D9, 16'hFE9C, 16'hD453, 16'hAC11, 16'hFEDD, 16'hF6DC, 16'hCCD5, 16'hD556, 16'hF69C, 16'hEE9C, 16'hEE9B, 16'hDD97, 16'hDD98, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hE65B, 16'hE61A, 16'hDE19, 16'hDE1A, 16'hDE19, 16'hDDD9, 16'hDDD8, 16'hDDD8, 16'hE69B, 16'hEE5B, 16'hDDD9, 16'hBC94, 16'hA411, 16'hBD15, 16'hDE1A, 16'hDE1A, 16'hDE1A, 16'hE61A, 16'hCD97, 16'h6A48, 16'h940F, 16'h8C10, 16'h8C0F, 16'h9450, 16'h9C92, 16'hA4D3, 16'hACD3, 16'h8BCF, 16'h93CF, 16'h8B8E, 16'hA4D3, 16'hAD14, 16'hAD14,
        16'hAD14, 16'hB514, 16'h8C0F, 16'hA4D3, 16'hCE18, 16'hC5D7, 16'hCE18, 16'hB555, 16'h9C92, 16'hFFDF, 16'hFFDF, 16'hAD14, 16'h94D2, 16'h83CF, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h4902, 16'hC596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h8490, 16'h84D0, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'h92CC, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hEE5A, 16'h8A8B, 16'hC596, 16'hFFDF, 16'hCDD7, 16'hCD56, 16'hCD57, 16'hA411, 16'hBD14, 16'hDE19, 16'hDE5A, 16'hDE5A, 16'hDE5A, 16'hDE59, 16'hB514, 16'hACD3, 16'hCDD8, 16'hD5D8, 16'hD5D8, 16'hCD97, 16'h728B, 16'h730C, 16'h7B0C, 16'h93CF, 16'hE619, 16'h7A8B, 16'hBD14, 16'hEE9B, 16'hE65A, 16'hEE9B,
        16'hE65A, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE61A, 16'hD557, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hC493, 16'hC3D1, 16'hF65A, 16'hFF1D, 16'hF6DC, 16'hF6DD, 16'hEE5A, 16'hA38F, 16'h6105, 16'h4904, 16'h3000, 16'h4104, 16'h3800, 16'h5000, 16'hCD15, 16'hFF1D, 16'hFF9F, 16'hFF5E, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1E, 16'hFEDD, 16'hFF1D, 16'hFE9C, 16'hFE9C, 16'hFF1D, 16'hF65C, 16'hFE9C, 16'hFEDD, 16'hF65B, 16'hF65C, 16'hFE9C, 16'hF61A, 16'hF61B, 16'hFE9D, 16'hF5DA, 16'hF61A, 16'hFE5C,
        16'hF5DA, 16'hF65B, 16'hF61A, 16'hED99, 16'hFE5B, 16'hF5D9, 16'h9A4B, 16'hE5D9, 16'hF6DD, 16'hEE5B, 16'hB411, 16'hE619, 16'hF69C, 16'hEE9C, 16'hEE5B, 16'hD557, 16'hE5D9, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hE65A, 16'hE619, 16'hDE1A, 16'hE61A, 16'hE619, 16'hDE19, 16'hDDD8, 16'hDDD9, 16'hE65A, 16'hE65A, 16'hDDD8, 16'hB452, 16'hAC11, 16'hBCD4, 16'hDE19, 16'hDE1A, 16'hDE1A, 16'hE61A, 16'hCD97, 16'h6A49, 16'h940F, 16'h8C50, 16'h8C0F, 16'h8C10, 16'h9C92, 16'hA4D3, 16'hA4D3, 16'h9410, 16'h8BCE, 16'h8B8E, 16'hACD3, 16'hAD14, 16'hAD14, 16'hAD14, 16'hB554, 16'h8C10, 16'hA492, 16'hCE18, 16'hC5D7, 16'hC618, 16'hC5D7, 16'h83CE, 16'hEF5D, 16'hFFDF, 16'hD659, 16'h8C91, 16'h7C0F, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'h8BCF, 16'h7B4C, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h7C4F, 16'h84D1, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE59, 16'h92CC, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hF71C, 16'hEE59, 16'h92CB, 16'hC555, 16'hFFDF, 16'hEF1D, 16'hB4D4, 16'hD597, 16'hAC52, 16'hAC93, 16'hD5D8, 16'hE65A, 16'hDE19, 16'hDE19, 16'hDE59, 16'hC597, 16'h9C51, 16'hBD15, 16'hCDD7, 16'hCDD8, 16'hD5D8, 16'hC556, 16'h9BD0, 16'h6A49, 16'h6A8A, 16'h8B4E, 16'hD598, 16'h6A09, 16'hCD56, 16'hE69B, 16'hE65A, 16'hEE9B, 16'hDE19, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5A, 16'hD557, 16'hE619, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hDD97, 16'hAACC, 16'hF619, 16'hFF1D, 16'hFF5E, 16'hF69B, 16'hAB8F, 16'h4000, 16'h48C4, 16'h3801, 16'h4104, 16'h1800, 16'h824A, 16'hE61A, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hFF1E,
        16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFEDD, 16'hFEDD, 16'hFEDD, 16'hFE9C, 16'hFF1D, 16'hFE9C, 16'hFE9C, 16'hFEDD, 16'hFE9C, 16'hF65B, 16'hFE9C, 16'hF65B, 16'hF61A, 16'hFEDD, 16'hF65B, 16'hF61A, 16'hFE5B, 16'hF61A, 16'hF65B, 16'hF61A, 16'hF5D9, 16'hF65B, 16'hF61B, 16'hDC95, 16'hA34E, 16'hF69B, 16'hF6DC, 16'hCD16, 16'hC493, 16'hEE9B, 16'hEE9B, 16'hF69C, 16'hEE5A, 16'hD557, 16'hE619, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE619, 16'hDE19, 16'hD5D8, 16'hDDD9, 16'hE65A, 16'hE65A, 16'hDDD8, 16'hA3D0, 16'hAC52, 16'hB4D4, 16'hDE59, 16'hDE5A, 16'hDE19, 16'hDE1A, 16'hCD56, 16'h6A08, 16'h940F,
        16'h8C50, 16'h8C0F, 16'h9450, 16'hA4D2, 16'hA492, 16'hA4D3, 16'h93D0, 16'h93CF, 16'h93CF, 16'hACD3, 16'hAD14, 16'hAD14, 16'hAD14, 16'hAD54, 16'h9451, 16'h9451, 16'hCE18, 16'hC5D7, 16'hC5D7, 16'hCE58, 16'h83CE, 16'hD69A, 16'hFFDF, 16'hEF5C, 16'h8C51, 16'h94D2, 16'h9C92, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD96, 16'h3000, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h7C4F, 16'h84D1, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69B, 16'h92CC, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hEE9B, 16'hEE5A, 16'h930D, 16'hB4D3, 16'hFFDF, 16'hFFDF, 16'hC596, 16'hCD56, 16'hC556, 16'hAC52, 16'hC556, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE5A, 16'hD619, 16'hAC93, 16'hA451, 16'hC556, 16'hCDD8, 16'hCDD7,
        16'hD5D8, 16'hB4D4, 16'h9C11, 16'h9C10, 16'h51C7, 16'h6A8A, 16'hCD16, 16'h6A09, 16'hD5D8, 16'hE65B, 16'hE65B, 16'hE69B, 16'hD5D8, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hDDD8, 16'hDD98, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE619, 16'h924A, 16'hE597, 16'hFF1D, 16'hFF5E, 16'hF61A, 16'hAB0E, 16'h3800, 16'h4001, 16'h4104, 16'h2800, 16'hA38F, 16'hFEDC, 16'hFF5F, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1D, 16'hFF1D, 16'hFEDD, 16'hFF1D, 16'hFEDD, 16'hFEDD, 16'hFEDD, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hEE5A, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFEDD, 16'hFF1E, 16'hF69D, 16'hFF1D, 16'hFEDD, 16'hF69C,
        16'hFEDD, 16'hFEDD, 16'hF65B, 16'hFE9C, 16'hFE9C, 16'hF61A, 16'hFE9C, 16'hFE9C, 16'hF61A, 16'hFE9C, 16'hF65B, 16'hF65B, 16'hFE5B, 16'hED99, 16'hFE5C, 16'hF61B, 16'hFE1A, 16'hB3D1, 16'hCD15, 16'hFEDD, 16'hEE5B, 16'hABD1, 16'hDD98, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5A, 16'hD597, 16'hE61A, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE61A, 16'hDE19, 16'hDE19, 16'hDDD8, 16'hDE19, 16'hE65A, 16'hE65A, 16'hD597, 16'h9B4E, 16'hAC52, 16'hB493, 16'hDE19, 16'hDE5A, 16'hDE19, 16'hE65A, 16'hCD56, 16'h6208, 16'h940F, 16'h8C10, 16'h8C0F, 16'h9450, 16'hA4D2, 16'h9C92, 16'hA4D3, 16'h8BCF, 16'h93CF, 16'h8B8E, 16'hA4D3, 16'hAD14, 16'hAD14, 16'hAD14, 16'hAD14, 16'h9451, 16'h9451, 16'hC617, 16'hC5D7, 16'hC5D7, 16'hD659, 16'h9491, 16'hBD95, 16'hFFDF, 16'hFFDF, 16'hA4D3, 16'h9512, 16'h7B8E, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h4904, 16'hA492, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C4F, 16'h8490, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h930D, 16'hEE9B, 16'hFFDF, 16'hFF9E, 16'hEEDC, 16'hE65A, 16'hEE19, 16'h934D, 16'h9C51, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hBCD4, 16'hDDD8, 16'hB493, 16'hBCD4, 16'hDDD8, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE59, 16'hBD56, 16'h9C51, 16'hAC93, 16'hC596, 16'hCDD7, 16'hCDD7, 16'hCD97, 16'hA492, 16'h9410, 16'hA492, 16'h93CF, 16'h3000, 16'h9BD0, 16'h8B0D, 16'hE61A, 16'hE65A, 16'hE65B, 16'hE65B, 16'hD598, 16'hE61A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hDDD9, 16'hD557, 16'hEE5B, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF69B, 16'hAB8F, 16'hCC94, 16'hFEDD, 16'hFF5E, 16'hCC94, 16'h1800, 16'h5000, 16'h824A, 16'h1000, 16'hB412, 16'hFEDD, 16'hFF1E, 16'hFF1D, 16'hFF1D, 16'hFEDD,
        16'hFEDD, 16'hFEDD, 16'hFEDD, 16'hFE9C, 16'hFEDD, 16'hF69C, 16'hFEDD, 16'hFEDC, 16'hFF1D, 16'hFEDD, 16'hFF1D, 16'hFEDD, 16'hFF1D, 16'hFF1E, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF1E, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF1D, 16'hFF1E, 16'hFF1D, 16'hFEDD, 16'hFF1E, 16'hFE9C, 16'hFEDD, 16'hFEDD, 16'hFE9C, 16'hFE9C, 16'hFEDD, 16'hF61B, 16'hFE9C, 16'hFEDD, 16'hF61A, 16'hFE5C, 16'hFE9C, 16'hFE5C, 16'hFE5C, 16'hF5D9, 16'hF65B, 16'hFE5C, 16'hF5D9, 16'hE598, 16'h9B0D, 16'hF65B, 16'hF6DC, 16'hCD15, 16'hBC12, 16'hEE5A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE619, 16'hD597, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE61A, 16'hDE19, 16'hDE19, 16'hD5D8, 16'hDE19, 16'hE65A,
        16'hE65B, 16'hCD56, 16'h8B0D, 16'hB493, 16'hAC52, 16'hD5D8, 16'hDE1A, 16'hDE19, 16'hDE5A, 16'hC556, 16'h6A08, 16'h9450, 16'h8C50, 16'h8C0F, 16'h9451, 16'hA4D3, 16'hA4D2, 16'hA4D3, 16'h8BCF, 16'h93CF, 16'h8B8E, 16'hAD13, 16'hAD14, 16'hAD14, 16'hAD14, 16'hAD14, 16'h9C92, 16'h9451, 16'hC617, 16'hC5D7, 16'hBDD7, 16'hCE59, 16'hAD55, 16'h9491, 16'hFFDF, 16'hFFDF, 16'hCE18, 16'h8CD2, 16'h7C4F, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h730C, 16'h730B, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD13, 16'h6B8D, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h9B4D, 16'hE69A, 16'hFFDF, 16'hF71C, 16'hE65A, 16'hE61A, 16'hE619, 16'h938F, 16'h8B8E, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hC556, 16'hD597, 16'hCD56, 16'hB4D3,
        16'hCD97, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE65A, 16'hD5D8, 16'h9C11, 16'h9C51, 16'hAC93, 16'hCD97, 16'hCDD7, 16'hD5D8, 16'hC556, 16'h9C51, 16'h9C11, 16'h9C51, 16'hA451, 16'h72CB, 16'h2800, 16'h6A49, 16'hDDD9, 16'hE65B, 16'hE65A, 16'hE65A, 16'hD597, 16'hDDD9, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE61A, 16'hE61A, 16'hD556, 16'hE619, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hF69C, 16'hCCD4, 16'h9ACD, 16'hFEDD, 16'hE5D9, 16'h6000, 16'h6146, 16'hDD98, 16'hA38F, 16'hB3D1, 16'hFEDD, 16'hFF1E, 16'hFEDD, 16'hFEDD, 16'hFE9C, 16'hFE9C, 16'hF69C, 16'hFEDD, 16'hF69C, 16'hFE9C, 16'hF69C, 16'hFEDC, 16'hF69C, 16'hFEDD, 16'hFF1D, 16'hFEDC, 16'hFEDD, 16'hFEDD, 16'hFF1E, 16'hFF1D, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1E, 16'hFF1D, 16'hFF1E, 16'hFEDD, 16'hFEDD, 16'hFF1D, 16'hFEDD, 16'hFE9C, 16'hFF1D, 16'hF69C, 16'hF65C, 16'hFEDD, 16'hF65C, 16'hFE5C, 16'hFEDC, 16'hFE9C, 16'hFE9C, 16'hF61A, 16'hF65B, 16'hFE9C, 16'hF5DA, 16'hFE1B, 16'hAB8F, 16'hCD15, 16'hFE9C, 16'hE61A, 16'hABD0, 16'hDD97, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hDDD9, 16'hDDD8, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE19, 16'hDE19, 16'hD5D8, 16'hDE19, 16'hE65A, 16'hE65B, 16'hC515, 16'h930D, 16'hB493, 16'hAC52, 16'hCD97, 16'hDE5A, 16'hDE19, 16'hDE1A, 16'hC515, 16'h6207, 16'h8C50, 16'h8C50, 16'h8C10, 16'h9C91, 16'hA4D3, 16'hA4D2, 16'hA4D3, 16'h8BCF, 16'h93CF, 16'h8B8E, 16'hAD13, 16'hAD14, 16'hAD14, 16'hA514, 16'hAD14, 16'h9C92, 16'h8C50, 16'hC5D7, 16'hC617, 16'hBDD7, 16'hCE59, 16'hBDD7, 16'h7BCE, 16'hF75D, 16'hFFDF, 16'hE6DC, 16'h8C91, 16'h8C91, 16'hA513, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h8BCF, 16'h4985, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h730C, 16'h9411, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'h92CC, 16'hD5D7, 16'hFFDF, 16'hEF1C, 16'hDE59, 16'hDE19, 16'hE619, 16'h9B8F, 16'h728A, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'hBCD4, 16'hD5D7, 16'hBCD4, 16'hC515, 16'hD619, 16'hDE19, 16'hDE19, 16'hDE5A, 16'hE65A, 16'hBD15, 16'h9410, 16'hA451, 16'hACD3, 16'hCDD7, 16'hCD97, 16'hD5D8, 16'hB514, 16'h9C51, 16'h9C51, 16'hA451, 16'hA492, 16'h834E, 16'h61C8, 16'h5986, 16'hCD57, 16'hE65B, 16'hE65B, 16'hE65A, 16'hD597, 16'hDDD8, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE61A, 16'hE61A, 16'hDD97, 16'hD557, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE619, 16'h9A8C, 16'hED98,
        16'hAA8C, 16'hB34F, 16'hF69C, 16'hEE1A, 16'hCC12, 16'hFEDD, 16'hFF1D, 16'hFEDD, 16'hFEDC, 16'hFE9C, 16'hF65B, 16'hFE9C, 16'hF65B, 16'hFEDC, 16'hF65B, 16'hFE9C, 16'hF65B, 16'hFEDC, 16'hF69C, 16'hFEDD, 16'hFEDC, 16'hFEDD, 16'hFEDD, 16'hFEDD, 16'hFF1E, 16'hFEDD, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1D, 16'hFF1E, 16'hFF1D, 16'hFEDD, 16'hFF1D, 16'hFEDD, 16'hF69C, 16'hFEDD, 16'hFE9C, 16'hF69C, 16'hFEDD, 16'hFEDC, 16'hFE9C, 16'hF65B, 16'hF65B, 16'hFE9D, 16'hF65B, 16'hFE1B, 16'hDD17, 16'hA34F, 16'hF69B, 16'hF69C, 16'hBC52, 16'hC493, 16'hE5D9, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hDDD8, 16'hE619, 16'hEE9B, 16'hE65B, 16'hEE5B, 16'hEE5B,
        16'hE65B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE19, 16'hDE19, 16'hD5D8, 16'hE61A, 16'hE65A, 16'hE65B, 16'hB492, 16'h8B0D, 16'hB493, 16'hAC52, 16'hCD57, 16'hDE5A, 16'hDE19, 16'hDE5A, 16'hBD15, 16'h6248, 16'h8C50, 16'h8C50, 16'h8C10, 16'h9CD2, 16'hA4D3, 16'h9C92, 16'hACD3, 16'h9410, 16'h8BCE, 16'h8B8E, 16'hAD14, 16'hA513, 16'hAD14, 16'hAD14, 16'hAD14, 16'h9CD2, 16'h8C10, 16'hBDD7, 16'hBE17, 16'hBE17, 16'hC658, 16'hCE59, 16'h7BCD, 16'hE6DB, 16'hFFDF, 16'hFF9E, 16'h9CD2, 16'h8CD2, 16'h840F, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA492, 16'h3902, 16'hB555, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE18, 16'h6A8A, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hA38F, 16'hCD55, 16'hFF9F, 16'hEEDB, 16'hDE19, 16'hDE19,
        16'hDE19, 16'hA411, 16'h4000, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD96, 16'hCD56, 16'hCD56, 16'hBD14, 16'hCD97, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE5A, 16'hD5D8, 16'h9410, 16'hA451, 16'hA451, 16'hB514, 16'hCDD7, 16'hCDD7, 16'hC596, 16'hAC93, 16'hA451, 16'h9C51, 16'h9C51, 16'hACD3, 16'h838E, 16'h7A8B, 16'h830D, 16'hE619, 16'hE65A, 16'hE65B, 16'hE61A, 16'hD597, 16'hD5D8, 16'hE619, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE619, 16'hE61A, 16'hE619, 16'hCD15, 16'hEE5A, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF69B, 16'hA34E, 16'hCC12, 16'hED98, 16'hFEDC, 16'hFF1D, 16'hE516, 16'hF61A, 16'hFF1D, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hF65B, 16'hF65C, 16'hF65B, 16'hFE9C, 16'hF69C, 16'hF65B, 16'hF65B, 16'hF69C, 16'hFE9C, 16'hFE9C, 16'hFEDD, 16'hFE9C, 16'hFEDD, 16'hFEDC, 16'hFF1D, 16'hFF1D, 16'hFEDD, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1D, 16'hFF1E, 16'hFEDD, 16'hFEDD, 16'hFEDD, 16'hFEDC, 16'hFEDD, 16'hFEDD, 16'hFEDD, 16'hFE9C, 16'hF65B, 16'hFE9D, 16'hFE5C, 16'hF61A, 16'hFE5C, 16'h9B4E, 16'hDD97, 16'hFEDC, 16'hE5D8, 16'h930D, 16'hDD97, 16'hE5D9, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hDDD8, 16'hE61A, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE19, 16'hDE19, 16'hD5D8, 16'hE61A, 16'hE65A, 16'hE65A, 16'h9BD0, 16'h9B8F, 16'hB4D4, 16'hAC52, 16'hC556, 16'hDE5A, 16'hDE19, 16'hDE1A, 16'hBCD4, 16'h6247, 16'h8C50, 16'h844F, 16'h8C50, 16'hA513, 16'hA513, 16'hA4D2, 16'hA4D3, 16'h8BCF, 16'h8B8E, 16'h838D, 16'hAD14, 16'hAD14, 16'hA4D3, 16'hA514, 16'hA514, 16'h9CD3, 16'h8C51, 16'hBDD7, 16'hC617, 16'hBE17, 16'hC618,
        16'hCE99, 16'h840F, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hB555, 16'h9512, 16'h738D, 16'hE71B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB554, 16'h4985, 16'h9C51, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD618, 16'hA452, 16'hE6DC, 16'hFF9E, 16'hAC11, 16'hB452, 16'hFF9F, 16'hEEDC, 16'hDE19, 16'hDE19, 16'hDE19, 16'hAC52, 16'h4000, 16'hBD15, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'hBCD4, 16'hDDD8, 16'hCD56, 16'hCD56, 16'hD5D8, 16'hDE19, 16'hDE19, 16'hDE5A, 16'hDE5A, 16'hB4D4, 16'h8BCF, 16'hA492, 16'h9C51, 16'hB514, 16'hCDD7, 16'hCDD7, 16'hBD55, 16'hA452, 16'hA492, 16'hA452, 16'h9C51, 16'hACD3, 16'h7B4D, 16'h5987, 16'h830D, 16'hE619, 16'hE65A, 16'hE65B, 16'hE619, 16'hD597, 16'hDDD8, 16'hDDD8, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE619,
        16'hE65A, 16'hEE5A, 16'hD516, 16'hDD98, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hE65B, 16'hF69C, 16'hC4D4, 16'hA34F, 16'hFEDD, 16'hF6DD, 16'hF69C, 16'hF61B, 16'hFEDC, 16'hF69B, 16'hFE9C, 16'hF65B, 16'hF65B, 16'hF65B, 16'hFE5B, 16'hF61A, 16'hFE9C, 16'hF65B, 16'hFE9C, 16'hF65B, 16'hFE9C, 16'hF65B, 16'hFEDC, 16'hFEDD, 16'hF69C, 16'hFEDD, 16'hF69C, 16'hFF1D, 16'hFEDD, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1D, 16'hFF1D, 16'hFEDD, 16'hFEDD, 16'hFEDD, 16'hFEDD, 16'hFE9C, 16'hFE9D, 16'hFE9C, 16'hF61B, 16'hFE9C, 16'hD516, 16'hAB90, 16'hF65B, 16'hFE9C, 16'h9B8F, 16'hB452,
        16'hE619, 16'hE61A, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hDDD8, 16'hE65A, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE61A, 16'hDE19, 16'hDDD9, 16'hD5D8, 16'hDE19, 16'hE65A, 16'hE619, 16'h934E, 16'h9BD0, 16'hB493, 16'hAC52, 16'hC556, 16'hDE5A, 16'hDE19, 16'hDE1A, 16'hB493, 16'h5A48, 16'h9450, 16'h8C50, 16'h8C50, 16'hA514, 16'hA4D3, 16'hA4D3, 16'hAD13, 16'h838E, 16'h8B8E, 16'h8BCF, 16'hAD14, 16'hA513, 16'hA513, 16'hA514, 16'hA514, 16'h9CD3, 16'h9491, 16'hBDD7, 16'hBDD7, 16'hBE17, 16'hBE17, 16'hCE99, 16'h8C90, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hC5D7, 16'h8CD1, 16'h73CD, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC5D7, 16'h5A48, 16'h838E, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hCDD7, 16'hA38F, 16'hAB90, 16'hFF5E, 16'hEF1C, 16'hD619, 16'hDE19, 16'hDE5A, 16'hAC93, 16'h6146, 16'h830C, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC556, 16'hCD57, 16'hD5D8, 16'hCD97, 16'hD597, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE65A, 16'hD5D8, 16'h8BCF, 16'h9C51, 16'hA492, 16'h9C51, 16'hB514, 16'hCD97, 16'hCD97, 16'hB4D4, 16'hA452, 16'hA492, 16'hA492, 16'hA492, 16'hACD3, 16'h834D, 16'h6A09, 16'h938E, 16'hE65A, 16'hE65A, 16'hE65B, 16'hDE19, 16'hD598, 16'hE61A, 16'hDDD8, 16'hE619, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hE619, 16'hE65A, 16'hEE5B, 16'hDDD8, 16'hC4D4, 16'hEE5B, 16'hEE5B, 16'hEE5A, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hE619, 16'h928B, 16'hEDD9, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE5B, 16'hFE5B, 16'hF61A, 16'hF61B, 16'hF61A, 16'hF65B, 16'hF61A, 16'hF65B, 16'hFE5C, 16'hF65B, 16'hFE5C, 16'hF65B, 16'hFE9C, 16'hF65B, 16'hFEDD, 16'hFE9C, 16'hFE9C, 16'hFEDD, 16'hFEDC, 16'hFF1D, 16'hFEDD, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F,
        16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFEDD, 16'hFEDD, 16'hFEDD, 16'hFE9C, 16'hF69C, 16'hFE5B, 16'h9B0D, 16'hE598, 16'hFE9C, 16'hD556, 16'h6145, 16'hE5D8, 16'hDDD9, 16'hE65A, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hE65A, 16'hDDD9, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD5D8, 16'hE65A, 16'hEE5B, 16'hDDD8, 16'h7A8A, 16'hA411, 16'hB493, 16'hAC52, 16'hBD15, 16'hDE5A, 16'hDE19, 16'hDE1A, 16'hAC52, 16'h5A47, 16'h9490, 16'h8C4F, 16'h9491, 16'hA513, 16'hA513, 16'hA4D3, 16'hA4D3, 16'h838E, 16'h8B8E,
        16'h8BCF, 16'hAD14, 16'hA513, 16'hA513, 16'hA514, 16'hA514, 16'h9CD3, 16'h8C51, 16'hBDD7, 16'hBE17, 16'hBE17, 16'hBE18, 16'hCE9A, 16'h9512, 16'hA513, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h8C91, 16'h844F, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h62CB, 16'h6ACB, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD618, 16'h928B, 16'hF6DC, 16'hF75D, 16'hD619, 16'hD619, 16'hDE5A, 16'hB514, 16'h938E, 16'h7A4A, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'hBCD4, 16'hDDD8, 16'hCD97, 16'hD5D7, 16'hD5D8, 16'hDE19, 16'hDE19, 16'hDE59, 16'hDE59, 16'hACD3, 16'h838E, 16'hA492, 16'h9C51, 16'h9C51, 16'hBD55, 16'hCD97, 16'hC596, 16'hAC93, 16'hA492, 16'hA492, 16'hA492, 16'hA492, 16'hACD3, 16'h830D, 16'h6A49, 16'h9BCF,
        16'hE65A, 16'hE65A, 16'hE65B, 16'hDE19, 16'hD598, 16'hEE5A, 16'hDE19, 16'hD5D8, 16'hEE5B, 16'hEE9C, 16'hEE9B, 16'hE619, 16'hE65A, 16'hE65B, 16'hE65A, 16'hC4D4, 16'hDD97, 16'hEE9B, 16'hE65A, 16'hE65A, 16'hEE5B, 16'hE65A, 16'hF69B, 16'hABD0, 16'hBC11, 16'hFE9C, 16'hFE5B, 16'hF61A, 16'hFE1A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF5DA, 16'hFE5B, 16'hF61A, 16'hFE9C, 16'hF65A, 16'hF65B, 16'hF65B, 16'hF69C, 16'hFE5B, 16'hFE9C, 16'hFEDD, 16'hFE9C, 16'hFEDC, 16'hFEDD, 16'hFEDD, 16'hFF1D, 16'hFEDD, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1D,
        16'hFF1D, 16'hFEDD, 16'hFEDD, 16'hFE9C, 16'hFEDD, 16'hC494, 16'hC493, 16'hFE9C, 16'hEDD9, 16'h7106, 16'h9B4E, 16'hE619, 16'hDDD8, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hE65A, 16'hDE19, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE19, 16'hDE19, 16'hDDD8, 16'hD5D8, 16'hE65A, 16'hE65B, 16'hCD56, 16'h6207, 16'hAC92, 16'hAC93, 16'hAC52, 16'hBD15, 16'hDE19, 16'hDE19, 16'hDE1A, 16'hAC12, 16'h6289, 16'h9491, 16'h8450, 16'h9CD2, 16'hA513, 16'hA4D3, 16'hA4D3, 16'hA4D3, 16'h834D, 16'h834D, 16'h8C10, 16'hA514, 16'hA514, 16'hA514, 16'h9D13, 16'hA514, 16'h9CD3, 16'h8C51, 16'hBE17, 16'hC617, 16'hBE17, 16'hBE17, 16'hCE9A, 16'h9D54, 16'h9491, 16'hFF9F, 16'hFFDF, 16'hE6DC, 16'h8C91, 16'h8490, 16'hAD14, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h734D, 16'h62CA, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h8A4B, 16'hE65A, 16'hFF9F, 16'hD619, 16'hD619, 16'hDE59, 16'hBD55, 16'h9BCF, 16'hA411, 16'hA452, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD96, 16'hD597, 16'hCD97, 16'hCDD7, 16'hCDD7, 16'hD619, 16'hDE19, 16'hDE19, 16'hDE59, 16'hCDD7, 16'h834E, 16'h9410, 16'h9C51, 16'h9C51, 16'h9C51, 16'hBD56, 16'hCD97, 16'hBD15, 16'hA492, 16'hAC93, 16'hA492, 16'hA493, 16'hACD3, 16'hACD4, 16'h834D, 16'h50C3, 16'hAC51, 16'hE65A, 16'hDE1A, 16'hE65A, 16'hDE19, 16'hD598, 16'hEE9B, 16'hDE19, 16'hDDD8, 16'hE61A, 16'hEE9C, 16'hEE9B, 16'hE619, 16'hE61A, 16'hE65A, 16'hE65A, 16'hDD98, 16'hB411, 16'hEE5B, 16'hEE5B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hDDD8, 16'h928A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF5D9, 16'hF65B, 16'hF61B, 16'hF65B, 16'hFE9C, 16'hF61A, 16'hFE9C, 16'hF65B, 16'hFE9C, 16'hF65B, 16'hFEDC, 16'hFEDD, 16'hFE9C,
        16'hFEDD, 16'hFE9C, 16'hFEDD, 16'hFEDD, 16'hFEDD, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFEDD, 16'hFF1E, 16'hEE1A, 16'hA38F, 16'hF61A, 16'hF65A, 16'h930D, 16'h920B, 16'hB452, 16'hE5D9, 16'hDDD9, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hE65A, 16'hE61A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE19, 16'hDE19, 16'hD5D8, 16'hD5D8, 16'hE65A, 16'hEE9B, 16'hB493, 16'h6248, 16'hAC93, 16'hAC93, 16'hAC92, 16'hBCD4, 16'hDE19, 16'hD619,
        16'hDE1A, 16'h9BD0, 16'h6ACA, 16'h9491, 16'h8C90, 16'hA513, 16'hA513, 16'hA513, 16'hA513, 16'hA4D2, 16'h7B4D, 16'h838E, 16'h9C92, 16'hA554, 16'hA514, 16'hA514, 16'h9D13, 16'hA514, 16'h9D13, 16'h8450, 16'hBDD7, 16'hBE17, 16'hBE17, 16'hBE18, 16'hCE9A, 16'hA5D5, 16'h8C90, 16'hF79E, 16'hFFDF, 16'hEF5D, 16'h94D1, 16'h8CD1, 16'h9C92, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDA, 16'h83CE, 16'h6B4B, 16'hC596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h9B8F, 16'hC515, 16'hFFDF, 16'hE69B, 16'hD619, 16'hDE59, 16'hCDD7, 16'h8B4E, 16'hC596, 16'h934F, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hC4D5, 16'hDDD8, 16'hCD97, 16'hD5D8, 16'hD5D8, 16'hDE19, 16'hDE19, 16'hD619, 16'hDE59, 16'hACD3, 16'h7B4D, 16'hA492, 16'h9C51, 16'h9C51, 16'hA452,
        16'hC556, 16'hC597, 16'hBD15, 16'hA493, 16'hA492, 16'hA492, 16'hA493, 16'hACD3, 16'hACD4, 16'h830D, 16'h7A4A, 16'hBCD3, 16'hEE5A, 16'hDE5A, 16'hE65A, 16'hDE19, 16'hD5D8, 16'hE65A, 16'hDE19, 16'hDDD8, 16'hDDD9, 16'hEE5B, 16'hEE9B, 16'hE619, 16'hE61A, 16'hE65A, 16'hE619, 16'hEE5A, 16'hA3D0, 16'hCD15, 16'hEE9B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hEE5B, 16'hA38E, 16'hD494, 16'hFE1A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF5DA, 16'hF5DA, 16'hF65B, 16'hF61A, 16'hFE9C, 16'hF65B, 16'hF65B, 16'hFE9C, 16'hF65B, 16'hFE9C, 16'hF65B, 16'hFEDC, 16'hFE9C, 16'hFE9C, 16'hFEDD, 16'hFE9C, 16'hFF1D, 16'hFEDD, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F,
        16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1D, 16'hFF1E, 16'hFEDD, 16'hB3D1, 16'hE598, 16'hFE9C, 16'h9B4F, 16'hB390, 16'hB390, 16'hC515, 16'hDDD8, 16'hE619, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE61A, 16'hE61A, 16'hDE19, 16'hDE19, 16'hD5D8, 16'hD5D8, 16'hDE5A, 16'hE65A, 16'h9B8F, 16'h72CB, 16'hACD3, 16'hAC93, 16'hAC92, 16'hB4D4, 16'hDE19, 16'hDE19, 16'hDE19, 16'h938F, 16'h734C, 16'h8C91, 16'h9491, 16'hA513, 16'hA513, 16'hA513, 16'hA514, 16'h9C51, 16'h730B, 16'h730B, 16'h9CD3, 16'h9D14, 16'h9D14, 16'h9D13, 16'h9D13, 16'hA554, 16'h9CD3, 16'h8450, 16'hBDD7, 16'hBE18, 16'hBE17, 16'hBE18, 16'hCE9A, 16'hADD6, 16'h8450, 16'hF75D, 16'hFFDF, 16'hF75E, 16'h9CD2, 16'h9512, 16'h9451, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h83CF,
        16'h734C, 16'hB555, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD15, 16'h9B4E, 16'hFF9E, 16'hEF1C, 16'hD618, 16'hD619, 16'hD619, 16'h938F, 16'hC556, 16'hC556, 16'hB492, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCDD8, 16'hCD56, 16'hCD97, 16'hD5D8, 16'hD618, 16'hD619, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD5D8, 16'h838E, 16'h8C10, 16'h9C92, 16'h9C51, 16'h9C51, 16'hA492, 16'hBD56, 16'hC597, 16'hB514, 16'hA493, 16'hA492, 16'hA492, 16'hA4D3, 16'hACD3, 16'hACD3, 16'h830D, 16'h6A08, 16'hBCD3, 16'hE65A, 16'hDE1A, 16'hE65A, 16'hDDD9, 16'hDDD8, 16'hDE19, 16'hDE19, 16'hDDD9, 16'hDDD8, 16'hE619, 16'hEE9B, 16'hDDD9, 16'hE619, 16'hEE5A, 16'hE619, 16'hEE5A, 16'hC515, 16'h7A09, 16'hE61A, 16'hEE5B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hD556, 16'hA28B, 16'hFE1A, 16'hF61A, 16'hF61A, 16'hF61A, 16'hF5DA, 16'hF65B,
        16'hF61B, 16'hF65B, 16'hFE9C, 16'hF61A, 16'hFE9C, 16'hF65B, 16'hFE9C, 16'hF69C, 16'hF69C, 16'hFEDD, 16'hFE9C, 16'hFE9C, 16'hFEDD, 16'hFEDD, 16'hFF1D, 16'hFEDD, 16'hFF1E, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1D, 16'hFF1E, 16'hC4D4, 16'hCC93, 16'hFE9C, 16'hBC53, 16'h928C, 16'hE556, 16'h8B0D, 16'hDDD8, 16'hDD98, 16'hE65A, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE61A, 16'hE61A, 16'hDE19, 16'hDE19,
        16'hD597, 16'hD5D9, 16'hE65A, 16'hE619, 16'h728A, 16'h838E, 16'hB4D3, 16'hAC92, 16'hAC92, 16'hB4D4, 16'hD619, 16'hDE19, 16'hDE19, 16'h834D, 16'h738D, 16'h9491, 16'h9CD2, 16'hA514, 16'hA513, 16'hA514, 16'hAD14, 16'h9410, 16'h730C, 16'h83CF, 16'hA514, 16'h9D13, 16'hA554, 16'hA514, 16'h9D13, 16'hA554, 16'h9D13, 16'h8450, 16'hBE17, 16'hBE18, 16'hBE18, 16'hBE58, 16'hCE9A, 16'hB658, 16'h94D1, 16'hEF5D, 16'hFFDF, 16'hFF9F, 16'hA513, 16'h94D2, 16'h9450, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h840F, 16'h7BCD, 16'hAD14, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h7A0A, 16'hE65A, 16'hF75D, 16'hD618, 16'hD618, 16'hD619, 16'hAC93, 16'hA451, 16'hEF1C, 16'h938F, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hC515, 16'hCD55, 16'hCD56, 16'hD619,
        16'hD619, 16'hDE19, 16'hDE19, 16'hD619, 16'hDE19, 16'hBD15, 16'h734C, 16'h9C92, 16'h9C51, 16'h9C51, 16'h9C51, 16'hA492, 16'hC556, 16'hC596, 16'hACD3, 16'hA492, 16'hA4D3, 16'hA492, 16'hA4D3, 16'hACD4, 16'hACD3, 16'h7ACB, 16'h6987, 16'hC515, 16'hE65A, 16'hDE5A, 16'hDE19, 16'hD5D8, 16'hDDD9, 16'hDE19, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hEE5B, 16'hE619, 16'hE619, 16'hEE5A, 16'hE619, 16'hE65A, 16'hDDD9, 16'h6987, 16'hAC51, 16'hF69C, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hEE5A, 16'h9ACD, 16'hDCD5, 16'hFE5B, 16'hF61A, 16'hF61A, 16'hF61A, 16'hFE5B, 16'hF61A, 16'hFE9C, 16'hFE5B, 16'hF61A, 16'hFE9C, 16'hF65B, 16'hFE9C, 16'hF69C, 16'hFEDD, 16'hFEDD, 16'hFE9C, 16'hFEDD, 16'hFEDD, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hF71D, 16'hF6DC, 16'hEE9B, 16'hEE5A, 16'hE619, 16'hE5D9, 16'hDD97,
        16'hDD97, 16'hDD97, 16'hE65A, 16'hF6DC, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1D, 16'hFF5E, 16'hDDD8, 16'hB38F, 16'hFE5B, 16'hC494, 16'h8209, 16'hF5D8, 16'hCC93, 16'hA3D0, 16'hE619, 16'hD598, 16'hE65A, 16'hE65B, 16'hEE5B, 16'hEE5B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE61A, 16'hDE1A, 16'hDE19, 16'hDE19, 16'hD597, 16'hDDD9, 16'hE65A, 16'hD597, 16'h51C5, 16'h8C10, 16'hACD3, 16'hAC93, 16'hAC92, 16'hB4D3, 16'hD5D8, 16'hDE19, 16'hD5D9, 16'h7ACC, 16'h7B8D, 16'h94D2, 16'hA513, 16'hA513, 16'hA513, 16'hA513, 16'hAD14, 16'h838E, 16'h6289, 16'h8C50, 16'hA554, 16'hA514, 16'hA513, 16'hA514, 16'h9D13, 16'hA554, 16'h94D2, 16'h8C51, 16'hBE17, 16'hBE18, 16'hBE18, 16'hC658, 16'hD6DA, 16'hBE58, 16'h8CD1, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hAD14, 16'h8CD1,
        16'h9450, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h840F, 16'h7C0E, 16'hACD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h8B4E, 16'hBCD4, 16'hF71D, 16'hDE59, 16'hD618, 16'hD619, 16'hC556, 16'h82CC, 16'hEF1C, 16'hCDD7, 16'hAC93, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69B, 16'hBCD4, 16'hC515, 16'hD5D8, 16'hD619, 16'hD619, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD618, 16'h8BCF, 16'h83CF, 16'h9C91, 16'h9451, 16'h9C91, 16'h9451, 16'hA493, 16'hC596, 16'hBD55, 16'hA493, 16'hACD3, 16'hA4D3, 16'hA4D3, 16'hACD3, 16'hACD4, 16'hACD3, 16'h7ACB, 16'h7208, 16'hC515, 16'hE65A, 16'hDE5A, 16'hCD97, 16'hD598, 16'hDE19, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hE61A, 16'hE619, 16'hE619, 16'hEE5A, 16'hE619, 16'hE61A, 16'hEE5A, 16'hABD1, 16'h6040, 16'hCD15,
        16'hF69B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hCCD4, 16'hA2CC, 16'hFE1A, 16'hF5DA, 16'hF61B, 16'hFE5C, 16'hF61A, 16'hF65B, 16'hFE9C, 16'hF65B, 16'hFE9C, 16'hFE9C, 16'hF69C, 16'hFEDC, 16'hF69C, 16'hFEDD, 16'hFF1D, 16'hFEDC, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFFDF, 16'hFF5E, 16'hEE9C, 16'hE61A, 16'hE61A, 16'hEE5A, 16'hEE9B, 16'hF69B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF69B, 16'hDD57, 16'hE65A, 16'hE619, 16'h9ACC, 16'h7003, 16'h830B, 16'hB4D3, 16'hDE5A, 16'hFF5E, 16'hFFDF, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF5F, 16'hE61A, 16'hBB4E, 16'hFDD9, 16'hC453, 16'h828B, 16'hE557, 16'hFE5B, 16'hA34E, 16'hC515, 16'hE619, 16'hDDD8, 16'hEE9B, 16'hEE5B, 16'hE65B, 16'hEE5B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A,
        16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE1A, 16'hDE19, 16'hDE19, 16'hDDD9, 16'hCD97, 16'hDE19, 16'hE65A, 16'hC515, 16'h49C5, 16'h9C91, 16'hB493, 16'hAC93, 16'hAC92, 16'hB493, 16'hD5D8, 16'hDE19, 16'hD598, 16'h6A8A, 16'h840F, 16'h9D13, 16'hA513, 16'h9D13, 16'hA513, 16'hA514, 16'hAD14, 16'h734D, 16'h6ACB, 16'h9CD3, 16'hA554, 16'h9D13, 16'hA513, 16'h9D13, 16'h9D13, 16'hA554, 16'h94D2, 16'h8C51, 16'hBE18, 16'hBE58, 16'hBE58, 16'hC659, 16'hD6DA, 16'hB657, 16'h8CD1, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hB555, 16'h8CD1, 16'h8C50, 16'hF79D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h840F, 16'h8450, 16'hA492, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC596, 16'h7A8B, 16'hE69A, 16'hDE9A, 16'hD618, 16'hCE18, 16'hCDD8, 16'h8B4D, 16'hCDD7,
        16'hFF9E, 16'h938E, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD5D7, 16'hBCD4, 16'hC515, 16'hD619, 16'hD619, 16'hDE19, 16'hDE19, 16'hD619, 16'hDE19, 16'hBD55, 16'h730C, 16'h9451, 16'h9C51, 16'h9C51, 16'h9C51, 16'h9450, 16'hA4D3, 16'hC596, 16'hB514, 16'hA493, 16'hACD3, 16'hA4D3, 16'hA492, 16'hACD3, 16'hACD4, 16'hA492, 16'h82CB, 16'h7A49, 16'hCD56, 16'hE65A, 16'hDE59, 16'hBCD4, 16'hD598, 16'hDE19, 16'hDDD9, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD9, 16'hE619, 16'hE619, 16'hDDD9, 16'hE65A, 16'hE61A, 16'hE619, 16'hEE5B, 16'hC4D5, 16'h92CB, 16'h828B, 16'hDDD8, 16'hEE9B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hEE1A, 16'h9ACC, 16'hD494, 16'hFE1B, 16'hF65B, 16'hFE5B, 16'hF65A, 16'hFE9C, 16'hFE9C, 16'hF65B, 16'hFEDD, 16'hF65B, 16'hFEDC, 16'hF6DC, 16'hFE9C, 16'hFF1D, 16'hFEDD, 16'hFEDC, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFFDF, 16'hFF1E, 16'hDE19,
        16'hDD97, 16'hE5D9, 16'hF6DC, 16'hFF5E, 16'hFF5E, 16'hFF1D, 16'hF69C, 16'hF65A, 16'hE5D8, 16'hE557, 16'hDCD4, 16'hCB90, 16'hE598, 16'hE619, 16'hC34F, 16'hD34F, 16'hBACD, 16'h7803, 16'h3000, 16'h7A8A, 16'hC556, 16'hFF5D, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hE65A, 16'hBB8F, 16'hF597, 16'hB3D0, 16'h8A8B, 16'hED58, 16'hFE9C, 16'hEE1A, 16'h8A4A, 16'hE5D8, 16'hDDD8, 16'hE619, 16'hEE5B, 16'hE65B, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE1A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE61A, 16'hDE19, 16'hDE19, 16'hDDD8, 16'hD598, 16'hDE19, 16'hE65A, 16'h9BCF, 16'h5248, 16'hA492, 16'hAC93, 16'hB493, 16'hAC93, 16'hAC93, 16'hCDD8, 16'hDE19, 16'hC556, 16'h51C7, 16'h9491, 16'h9D13, 16'h9D13, 16'h9D13, 16'hA514, 16'hAD54, 16'hA4D3, 16'h628A, 16'h6B0C, 16'hA514, 16'hA554, 16'hA514, 16'h9D14, 16'h9D14, 16'h9D14, 16'hAD55, 16'h94D2, 16'h8C51,
        16'hBE18, 16'hBE18, 16'hBE58, 16'hC699, 16'hD6DB, 16'hB658, 16'h94D2, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8490, 16'h9450, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE17, 16'h8C50, 16'h8450, 16'hA4D3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h728B, 16'hB514, 16'hE69A, 16'hD659, 16'hD618, 16'hD659, 16'h9C51, 16'hA411, 16'hFFDF, 16'hCDD7, 16'hAC52, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hC515, 16'hB452, 16'hCD97, 16'hDE19, 16'hD619, 16'hD619, 16'hD619, 16'hD619, 16'hD619, 16'h9C11, 16'h7B8D, 16'h9C91, 16'h9C91, 16'h9C91, 16'h9451, 16'h9450, 16'hACD3, 16'hBD96, 16'hACD4, 16'hACD3, 16'hA4D3, 16'hA4D3, 16'hA493, 16'hA4D3, 16'hAD14, 16'h9C92, 16'h82CB, 16'h7A4A, 16'hCD56, 16'hDE5A, 16'hDE19, 16'hA411, 16'hD598, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19,
        16'hDE19, 16'hDE19, 16'hE619, 16'hE619, 16'hDDD9, 16'hE61A, 16'hE61A, 16'hE619, 16'hE61A, 16'hD597, 16'h8B0C, 16'hAC52, 16'h6A09, 16'hD597, 16'hEE9B, 16'hDE19, 16'hE61A, 16'hEE5B, 16'hCD15, 16'h9ACC, 16'hFE1A, 16'hFE9C, 16'hF65B, 16'hFE9C, 16'hFE9C, 16'hF69B, 16'hFE9C, 16'hFEDC, 16'hF69C, 16'hFEDD, 16'hFEDD, 16'hFEDD, 16'hFF1D, 16'hFEDD, 16'hFEDD, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF5F, 16'hD5D8, 16'hCD15, 16'hE619, 16'hF71D, 16'hF6DC, 16'hF65B, 16'hE557, 16'hDC93, 16'hCB90, 16'hCB0F, 16'hCACE, 16'hCA8D, 16'hCA8E, 16'hD2CE, 16'hD30F, 16'hCA8D, 16'hC24C, 16'hD350, 16'hD350, 16'hDB91, 16'hD3D1, 16'hBB0E, 16'h78C5, 16'h000, 16'h7208, 16'hE69A, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hEE5A, 16'hC411, 16'hDC94, 16'h9A8C, 16'hAB8F, 16'hF598, 16'hF61A, 16'hFF5F, 16'hCD56,
        16'h9B4E, 16'hE619, 16'hDDD8, 16'hE65A, 16'hEE5B, 16'hE65A, 16'hEE5B, 16'hE619, 16'hE619, 16'hE65A, 16'hE65A, 16'hDE19, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD5D8, 16'hD5D8, 16'hE65A, 16'hDDD9, 16'h61C7, 16'h634B, 16'hACD3, 16'hAC93, 16'hAC93, 16'hAC93, 16'hAC93, 16'hCDD8, 16'hDE5A, 16'hBCD4, 16'h5207, 16'h9CD3, 16'h9D13, 16'hA513, 16'hA513, 16'hA554, 16'hB555, 16'h8C10, 16'h59C7, 16'h7C0F, 16'hA554, 16'h9D14, 16'h9D14, 16'h9D14, 16'hA554, 16'h9D54, 16'hAD54, 16'h94D2, 16'h8C91, 16'hBE18, 16'hBE58, 16'hBE58, 16'hCE9A, 16'hDF1B, 16'hB618, 16'h94D2, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hAD54, 16'h7C4F, 16'h9491, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD95, 16'h8CD1, 16'h8491, 16'hAD14, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hACD3, 16'h6A8A, 16'hCE18, 16'hD659, 16'hCE18, 16'hD659, 16'hBD96, 16'h82CC, 16'hEEDB, 16'hFFDF, 16'h9410, 16'hD619, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'h9BD0, 16'hAC92, 16'hD619, 16'hD619, 16'hD619, 16'hD619, 16'hD619, 16'hD619, 16'hCD97, 16'h7B8D, 16'h8450, 16'h9C91, 16'h9C92, 16'h9491, 16'h9451, 16'h9450, 16'hAD14, 16'hBD55, 16'hACD3, 16'hACD3, 16'hA4D3, 16'hA4D3, 16'hA4D3, 16'hACD4, 16'hAD14, 16'h9C92, 16'h82CB, 16'h7A4A, 16'hD597, 16'hE65A, 16'hD618, 16'h8B4E, 16'hD598, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE619, 16'hE619, 16'hDDD9, 16'hE619, 16'hE61A, 16'hDDD9, 16'hDDD9, 16'hE61A, 16'h934E, 16'hB452, 16'hAC52, 16'h61C7, 16'hCD56, 16'hEE5A, 16'hDE19, 16'hDE19, 16'hEE5B, 16'hA34E, 16'hCCD4, 16'hFE9C, 16'hF65B, 16'hFE9C, 16'hFE9C, 16'hF69B, 16'hFEDD, 16'hFE9C, 16'hFE9C, 16'hFEDD, 16'hFEDD, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F,
        16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hEE5B, 16'h934E, 16'h5000, 16'hC4D4, 16'hFEDD, 16'hD4D4, 16'hCACE, 16'hD30F, 16'hCACD, 16'hD30F, 16'hD34F, 16'hD350, 16'hD350, 16'hD390, 16'hD350, 16'hD350, 16'hD350, 16'hD350, 16'hD390, 16'hD34F, 16'hD34F, 16'hCB4F, 16'hCB4F, 16'hD390, 16'hD390, 16'hAA8C, 16'h4800, 16'h4000, 16'hDE18, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hE619, 16'hBB0E, 16'hBB4F, 16'hAB0E, 16'hD494, 16'hFDD9, 16'hF65B, 16'hFF5E, 16'hFF5E, 16'hA3D0, 16'hC4D4, 16'hE619, 16'hDDD9, 16'hE65A, 16'hEE5B, 16'hE65A, 16'hEE5B, 16'hD597, 16'hDE19, 16'hE65A, 16'hDE19, 16'hDE19, 16'hDE1A, 16'hE61A, 16'hE61A, 16'hDE1A, 16'hE61A, 16'hE61A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD598, 16'hD5D8, 16'hEE5B, 16'hBCD5, 16'h3000, 16'h7BCE, 16'hB514, 16'hAC93, 16'hAC93, 16'hB4D3, 16'hAC92, 16'hCDD8, 16'hDE5A, 16'hAC52, 16'h62CA, 16'hA514, 16'h9D13, 16'hA514, 16'hA514, 16'hA554, 16'hA514,
        16'h6ACB, 16'h41C6, 16'h8C91, 16'hA554, 16'h9D14, 16'hA554, 16'h9D54, 16'hA554, 16'h9D54, 16'hA595, 16'h8C91, 16'h8C91, 16'hBE58, 16'hBE58, 16'hBE58, 16'hD6DB, 16'hDF1C, 16'hADD6, 16'h9CD2, 16'hF79E, 16'hFFDF, 16'hFF9F, 16'hA554, 16'h740E, 16'hA4D2, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h9C92, 16'h9553, 16'h8490, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'h5A07, 16'hA492, 16'hD659, 16'hCE18, 16'hCE18, 16'hCE59, 16'h8BCF, 16'hBD15, 16'hFFDF, 16'hE6DB, 16'h8B4E, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCDD7, 16'h828B, 16'hC556, 16'hDE59, 16'hD619, 16'hD619, 16'hD619, 16'hD619, 16'hD659, 16'hB4D4, 16'h6B4C, 16'h9491, 16'h9491, 16'h9491, 16'h9451, 16'h9451, 16'h9451, 16'hAD14, 16'hB555, 16'hA4D3, 16'hA4D3, 16'hA4D3, 16'hA4D3, 16'hA4D3, 16'hAD14, 16'hAD14,
        16'h9451, 16'h8B4D, 16'h828B, 16'hCD56, 16'hE65A, 16'hCD97, 16'h7A8B, 16'hD597, 16'hE61A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE619, 16'hE619, 16'hDE19, 16'hDDD9, 16'hE619, 16'hDDD9, 16'hDDD8, 16'hEE5B, 16'hB493, 16'hA3D0, 16'hCD56, 16'hA411, 16'h6145, 16'hBCD3, 16'hEE1A, 16'hE619, 16'hE65A, 16'hDD97, 16'h928A, 16'hF5D9, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFEDD, 16'hFEDC, 16'hFEDD, 16'hFF1D, 16'hFEDD, 16'hFF1E, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hCD56, 16'h6000, 16'h6000, 16'h8146, 16'hBA4B, 16'hCB0F, 16'hD30F, 16'hD350, 16'hD350, 16'hD350, 16'hD350, 16'hD350, 16'hD350, 16'hD350, 16'hD350, 16'hD350, 16'hD350, 16'hD350, 16'hD34F, 16'hD34F, 16'hCB4F, 16'hD34F, 16'hD34F, 16'hD34F, 16'hCB0F, 16'hCB4F, 16'hD350, 16'hBACD, 16'h5800, 16'h4800, 16'hEEDB, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF1E, 16'hC4D4, 16'h9106, 16'hB30E, 16'hD494, 16'hF599, 16'hF5D9, 16'hF65B, 16'hFF5E, 16'hFF9F, 16'hF69C, 16'h8A8C, 16'hD597, 16'hDDD9, 16'hDE19, 16'hE65A, 16'hE65B, 16'hE65B, 16'hE619, 16'hCD15, 16'hE65A, 16'hE65A, 16'hDE19, 16'hDE19, 16'hE65A, 16'hDE19, 16'hE619, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD598, 16'hDE19, 16'hEE5A, 16'h9BCF, 16'h3140, 16'h8C50, 16'hB514, 16'hACD3, 16'hB4D4, 16'hB493, 16'hAC52, 16'hCDD8, 16'hDE5A, 16'h8B4E, 16'h734C, 16'hA555, 16'hA514, 16'hA554, 16'hA513, 16'hA554, 16'h9491, 16'h4946, 16'h738D, 16'h94D2, 16'hA555, 16'hA554, 16'hA554, 16'hA554, 16'hA554, 16'h9D54, 16'hA595, 16'h8C91, 16'h9492, 16'hBE58, 16'hBE58, 16'hBE98, 16'hDF1B, 16'hE75C, 16'hAD95, 16'hA513, 16'hF79E, 16'hFFDF, 16'hF79E, 16'hA513, 16'h6B8C, 16'hB595, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h83CE, 16'hA595, 16'h740E, 16'hD658, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA492, 16'h49C6, 16'hBD97, 16'hD659, 16'hCE58, 16'hCE59, 16'hB555, 16'h8B4E, 16'hF75D, 16'hFFDF, 16'hC596, 16'hB4D4, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAC92, 16'h8B8E, 16'hD619, 16'hD619, 16'hD619, 16'hD619, 16'hD619, 16'hD619, 16'hD619, 16'h9410, 16'h73CE, 16'h94D2, 16'h9491, 16'h9491, 16'h9491, 16'h9491, 16'h9491, 16'hA514, 16'hAD54, 16'hAD13, 16'hAD13, 16'hA4D3, 16'hA4D3, 16'hA4D3, 16'hAD14, 16'hAD14, 16'h9492, 16'h934D, 16'h8ACC, 16'hD597, 16'hE65A, 16'hC556, 16'h6A09, 16'hD597, 16'hE65A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE619, 16'hE619, 16'hE619, 16'hE619, 16'hDDD9, 16'hDE19, 16'hDDD9, 16'hD598, 16'hEE5B, 16'hCD56, 16'hA38F, 16'hC515, 16'hCD56, 16'h934D, 16'h5000, 16'h9B8F, 16'hDD98, 16'hE61A, 16'hEE5A, 16'hCC94, 16'h9ACC, 16'hF65B, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFEDD, 16'hFEDD, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E,
        16'hFF1E, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hC515, 16'h3000, 16'h7105, 16'h7905, 16'hBA8C, 16'hDB50, 16'hD30F, 16'hD350, 16'hD34F, 16'hD34F, 16'hD34F, 16'hD350, 16'hD350, 16'hD350, 16'hD350, 16'hD34F, 16'hD34F, 16'hD34F, 16'hD34F, 16'hD34F, 16'hD34F, 16'hCB4F, 16'hCB0F, 16'hCB4F, 16'hCB4F, 16'hCB4F, 16'hCB4F, 16'hCB0F, 16'hD350, 16'hBACD, 16'h3800, 16'h938E, 16'hFF9F, 16'hFF5E, 16'hFF1E, 16'hF71D, 16'hF6DD, 16'hEE5B, 16'hD556, 16'hB38F, 16'hB390, 16'hE517, 16'hF5D9, 16'hFE1A, 16'hF61A, 16'hF6DC, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hD598, 16'h9B8F, 16'hE619, 16'hDDD9, 16'hDE19, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hC493, 16'hC4D4, 16'hEE5B, 16'hE61A, 16'hDDD9, 16'hDE19, 16'hDE19, 16'hDE1A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD9, 16'hCD97, 16'hE65A, 16'hDDD8, 16'h69C8, 16'h5247, 16'h9C92, 16'hB514, 16'hB4D4, 16'hB4D4,
        16'hACD3, 16'hA452, 16'hD618, 16'hD619, 16'h7ACC, 16'h840F, 16'hA554, 16'h9D14, 16'hA554, 16'hA554, 16'hA514, 16'h6ACB, 16'h5249, 16'h740F, 16'h9553, 16'hA554, 16'h9D54, 16'h9D54, 16'hA554, 16'hA554, 16'h9D54, 16'hA555, 16'h8C91, 16'h94D2, 16'hBE58, 16'hBE58, 16'hBE98, 16'hE75C, 16'hEF5D, 16'h9D13, 16'hAD54, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h9491, 16'h5288, 16'hCE58, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE18, 16'h7C4F, 16'hA5D5, 16'h7BCE, 16'hE71B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h4985, 16'h7B8E, 16'hCE18, 16'hCE59, 16'hCE58, 16'hCE19, 16'h8B8F, 16'hC596, 16'hFFDF, 16'hFFDE, 16'h9C50, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h830D, 16'hACD3, 16'hD659, 16'hD618, 16'hD619, 16'hD619, 16'hD619, 16'hD659, 16'hC597, 16'h6B0C, 16'h8490, 16'h94D2, 16'h9491, 16'h8C91,
        16'h8C91, 16'h9491, 16'h9491, 16'hA513, 16'hAD14, 16'hA513, 16'hAD14, 16'hA513, 16'hA4D3, 16'h9CD3, 16'hA514, 16'hAD14, 16'h9C92, 16'h8B0C, 16'h828B, 16'hCD56, 16'hDE5A, 16'hC556, 16'h61C8, 16'hCD96, 16'hE65A, 16'hDE1A, 16'hDE1A, 16'hDE1A, 16'hDE1A, 16'hDE19, 16'hDE19, 16'hE619, 16'hE619, 16'hDDD9, 16'hDDD9, 16'hDE19, 16'hCD57, 16'hE61A, 16'hDDD8, 16'hA3D0, 16'hC556, 16'hCD56, 16'h7A49, 16'hC411, 16'hAB8F, 16'h71C8, 16'hBC52, 16'hDD57, 16'hEDD8, 16'hB3D0, 16'hBC12, 16'hFE9D, 16'hFEDD, 16'hFEDD, 16'hFF1E, 16'hFEDD, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hD619, 16'h2800, 16'h6946, 16'h7083, 16'hB28C, 16'hD34F, 16'hCB4F, 16'hD34F, 16'hD34F, 16'hD34F, 16'hD34F, 16'hD350, 16'hD34F, 16'hD34F, 16'hD34F, 16'hD391, 16'hDBD2, 16'hE413, 16'hE453, 16'hE453, 16'hE454, 16'hE413, 16'hDBD2, 16'hD391, 16'hD390, 16'hCB0F, 16'hCB0E, 16'hCB0F,
        16'hCB4F, 16'hCB4F, 16'hDB50, 16'hB2CC, 16'h1800, 16'hD5D8, 16'hFF9F, 16'hF69C, 16'hE598, 16'hD515, 16'hD4D4, 16'hDD16, 16'hF5D9, 16'hFE5B, 16'hFE1B, 16'hF61B, 16'hF69C, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hB411, 16'hC515, 16'hE61A, 16'hDE19, 16'hE65A, 16'hE65A, 16'hE65B, 16'hE619, 16'h92CC, 16'hD597, 16'hE65A, 16'hDE19, 16'hD5D8, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD5D8, 16'hCD97, 16'hE61A, 16'hB453, 16'h5207, 16'h6B4B, 16'hA4D3, 16'hB514, 16'hB4D4, 16'hB4D4, 16'hAC93, 16'h9C11, 16'hD619, 16'hD5D8, 16'h6249, 16'h9CD2, 16'hA554, 16'h9D54, 16'h9D14, 16'hA554, 16'h9450, 16'h5248, 16'h73CE, 16'h744F, 16'h9D54, 16'hA554, 16'hA554, 16'h9D54, 16'hA554, 16'h9D54, 16'h9D54, 16'hA554, 16'h8C50, 16'h9CD3, 16'hBE58, 16'hBE98, 16'hBE59, 16'hEF5D, 16'hEF5D, 16'h8C50, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h7B8E, 16'h62CA, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFF9F, 16'h9C92, 16'h9593, 16'h9D54, 16'h9491, 16'hFFDE, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h9C51, 16'h6A8A, 16'hA4D2, 16'hCE59, 16'hCE59, 16'hCE59, 16'hB515, 16'h93CF, 16'hF75D, 16'hFFDF, 16'hEF1C, 16'h8BCF, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h724A, 16'hCD97, 16'hD659, 16'hD619, 16'hD619, 16'hD619, 16'hD618, 16'hD619, 16'hA492, 16'h5B0A, 16'h8CD2, 16'h94D2, 16'h8C91, 16'h8C91, 16'h8C91, 16'h8C91, 16'h9491, 16'hA514, 16'hA514, 16'hA514, 16'hA513, 16'hA513, 16'h9CD2, 16'h9CD3, 16'hA514, 16'hAD55, 16'h9491, 16'h930D, 16'h930C, 16'hD597, 16'hE65A, 16'hBD15, 16'h5987, 16'hC556, 16'hE65A, 16'hDE1A, 16'hDE1A, 16'hDE1A, 16'hDE1A, 16'hDE1A, 16'hDE19, 16'hE619, 16'hE61A, 16'hDE19, 16'hDDD9, 16'hDDD9, 16'hCD56, 16'hDE19, 16'hDE19, 16'hA3D0, 16'hCD56, 16'hBCD4, 16'h8208, 16'hCC94, 16'hCC94, 16'hAB4E, 16'h7042, 16'h8A8B,
        16'h92CC, 16'hC452, 16'hA28B, 16'hBC11, 16'hF61A, 16'hF65B, 16'hEDD9, 16'hF65B, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF1E, 16'h6A49, 16'h5800, 16'h68C4, 16'hA24A, 16'hD350, 16'hCB4F, 16'hD34F, 16'hD34F, 16'hD34F, 16'hD34F, 16'hD350, 16'hD34F, 16'hCB4F, 16'hDBD1, 16'hE454, 16'hEC95, 16'hECD5, 16'hF4D6, 16'hF4D6, 16'hECD6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hEC95, 16'hEC95, 16'hEC54, 16'hDC12, 16'hD390, 16'hCB4F, 16'hCB0F, 16'hCB4F, 16'hDB90, 16'h8084, 16'h934E, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hFEDD, 16'hFEDC, 16'hF6DC, 16'hFEDD, 16'hFF5F, 16'hFF9F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hF6DD, 16'h9B8F, 16'hE619, 16'hE619, 16'hDE19, 16'hE65A, 16'hE65A, 16'hEE5B, 16'hB411, 16'h930D, 16'hE61A, 16'hE65A, 16'hDDD9, 16'hD5D8, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19,
        16'hDE19, 16'hDDD9, 16'hCD97, 16'hD5D8, 16'hDDD8, 16'h7ACC, 16'h630B, 16'h734C, 16'hB514, 16'hB514, 16'hB514, 16'hB4D4, 16'hA452, 16'h9C11, 16'hDE59, 16'hC556, 16'h5207, 16'h9D13, 16'hA514, 16'hA554, 16'hA554, 16'h9D13, 16'h5A48, 16'h840F, 16'h744F, 16'h7C90, 16'h9D54, 16'hA595, 16'hA595, 16'hA554, 16'hA554, 16'h9D54, 16'hA595, 16'h9D14, 16'h7BCE, 16'h9D13, 16'hBE99, 16'hB698, 16'hC699, 16'hF79E, 16'hEF5D, 16'h7BCE, 16'hCE58, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h5207, 16'h9CD2, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h73CD, 16'hAE57, 16'h844F, 16'hCE17, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD658, 16'h838E, 16'h9C51, 16'hA4D3, 16'hCE59, 16'hCE59, 16'hCE18, 16'h8BCF, 16'hCDD7, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h9C51, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD55, 16'h834E, 16'hD619,
        16'hD619, 16'hD619, 16'hD619, 16'hD619, 16'hD619, 16'hCDD7, 16'h838E, 16'h7C0E, 16'h94D2, 16'h94D2, 16'h8C91, 16'h8C91, 16'h8C91, 16'h8C91, 16'h94D2, 16'hA514, 16'hAD54, 16'hA514, 16'hA514, 16'hA514, 16'h9491, 16'h9CD3, 16'hA554, 16'hAD55, 16'h9491, 16'h9B8E, 16'h930C, 16'hCD96, 16'hDE59, 16'hBD55, 16'h5145, 16'hBD15, 16'hE65A, 16'hDE19, 16'hDE1A, 16'hDE19, 16'hDE1A, 16'hDE1A, 16'hE619, 16'hE61A, 16'hE61A, 16'hDE19, 16'hDDD9, 16'hDDD9, 16'hCD56, 16'hDDD8, 16'hE61A, 16'hB493, 16'hCD16, 16'hAC11, 16'h9ACB, 16'hD4D5, 16'hC453, 16'hC411, 16'h9A4A, 16'hD4D4, 16'hDD16, 16'hBC52, 16'hC412, 16'hAACC, 16'hC3D1, 16'hE517, 16'hEE1A, 16'hFF1E, 16'hFF5E, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hCD97, 16'h2800, 16'h6945, 16'h8988, 16'hCB4F, 16'hCB4F, 16'hCB4F, 16'hD34F, 16'hD34F, 16'hCB4F, 16'hD34F, 16'hCB4F, 16'hD391, 16'hE454, 16'hECD6, 16'hF4D6, 16'hECD5,
        16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hECD5, 16'hEC95, 16'hEC95, 16'hECD5, 16'hF4D6, 16'hF4D5, 16'hEC95, 16'hEC54, 16'hDB91, 16'hCB0F, 16'hD350, 16'hCB0E, 16'h6002, 16'hEEDC, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF9F, 16'hD597, 16'hA411, 16'hEE5A, 16'hDE19, 16'hE61A, 16'hE65A, 16'hEE5B, 16'hDD98, 16'h70C4, 16'hB452, 16'hE65A, 16'hE61A, 16'hD5D8, 16'hDDD9, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD9, 16'hDE19, 16'hD598, 16'hCD97, 16'hDDD9, 16'hBCD4, 16'h5A49, 16'h738D, 16'h838E, 16'hBD55, 16'hB514, 16'hB4D4, 16'hBD15, 16'hA451, 16'hA492, 16'hDE5A, 16'hA452, 16'h5A89, 16'hA554, 16'hA514, 16'hA554, 16'hA513, 16'h62CA, 16'h840F, 16'h94D3, 16'h63CE, 16'h84D1, 16'hA595, 16'hA554, 16'h9D54, 16'hA554, 16'hA554, 16'hA554, 16'hA595, 16'h94D3, 16'h840F, 16'hA553, 16'hBE99, 16'hBE99, 16'hCE9A, 16'hFFDF, 16'hE71B, 16'h734C, 16'hE6DB, 16'hFFDF,
        16'hFFDF, 16'hC617, 16'h3900, 16'hD699, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h8C10, 16'h9553, 16'hA594, 16'h840F, 16'hF79D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h9C91, 16'hCDD7, 16'hB555, 16'hA4D3, 16'hCE59, 16'hD69A, 16'hB555, 16'h8B4D, 16'hEF1D, 16'hFFDF, 16'hFFDF, 16'hBD96, 16'hB514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h9410, 16'hA492, 16'hD659, 16'hD619, 16'hD618, 16'hD618, 16'hD618, 16'hD619, 16'hB4D4, 16'h9410, 16'h8450, 16'h94D2, 16'h94D2, 16'h8CD2, 16'h8CD2, 16'h8CD2, 16'h8C91, 16'h94D2, 16'hAD54, 16'hAD54, 16'hA514, 16'hA514, 16'hA514, 16'h9491, 16'h9D13, 16'hA554, 16'hA555, 16'h9C92, 16'h934D, 16'h82CB, 16'hCD56, 16'hDE59, 16'hB514, 16'h5185, 16'hB4D3, 16'hE65A, 16'hDE19, 16'hDE1A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE619, 16'hE61A, 16'hE619, 16'hDE19, 16'hDDD9,
        16'hCD56, 16'hCD57, 16'hEE5B, 16'hCD15, 16'hC4D4, 16'h92CB, 16'hB3CF, 16'hD4D4, 16'hCC93, 16'hCC53, 16'hA28B, 16'hBB8F, 16'hF5D9, 16'hFE1A, 16'hFE1A, 16'hFDD9, 16'hFE5B, 16'hFF5E, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'h93D0, 16'h4800, 16'h6904, 16'hB2CD, 16'hD350, 16'hCB4F, 16'hCB4F, 16'hD34F, 16'hD34F, 16'hCB4F, 16'hCB4F, 16'hDC13, 16'hECD5, 16'hECD6, 16'hEC95, 16'hEC95, 16'hECD5, 16'hF4D6, 16'hEC95, 16'hEC95, 16'hEC95, 16'hECD5, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hF495, 16'hE454, 16'hD390, 16'hDB90, 16'h8805, 16'hD619, 16'hFFDF, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5F, 16'hA410, 16'hC516, 16'hEE5A, 16'hE619, 16'hE61A, 16'hE65A, 16'hEE5A, 16'hA38E, 16'h7945, 16'hCD15, 16'hE65A,
        16'hDE19, 16'hD5D8, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD9, 16'hDE19, 16'hDDD8, 16'hCD56, 16'hD597, 16'hDDD8, 16'h834D, 16'h6B8D, 16'h630B, 16'h9C11, 16'hBD55, 16'hB515, 16'hB514, 16'hBD15, 16'h93CF, 16'hB4D4, 16'hDE59, 16'h8B4E, 16'h738D, 16'hA554, 16'hAD95, 16'hA554, 16'h6B0B, 16'h8C51, 16'hAD96, 16'h8C91, 16'h63CD, 16'h84D2, 16'hA595, 16'hA554, 16'hA595, 16'hA595, 16'hA554, 16'hA554, 16'hA595, 16'h8C91, 16'hA513, 16'hA595, 16'hBED9, 16'hBE98, 16'hDF1B, 16'hFFDF, 16'hD659, 16'h7B8D, 16'hF79D, 16'hFFDF, 16'hFFDF, 16'h9450, 16'h83CE, 16'hFFDE, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD96, 16'h740E, 16'hAE16, 16'h6B4C, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'hACD3, 16'hF79E, 16'hB555, 16'hA4D3, 16'hD69A, 16'hD69A, 16'h9451, 16'hB4D3, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hACD2, 16'hC5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'h7B0C, 16'hC556, 16'hD619, 16'hD618, 16'hD619, 16'hD619, 16'hD619, 16'hCDD8, 16'hA452, 16'hB555, 16'h73CF, 16'h9D13, 16'h9512, 16'h8CD1, 16'h8CD1, 16'h8C91, 16'h8C91, 16'h9CD2, 16'hAD55, 16'hA554, 16'hA514, 16'hA514, 16'hA514, 16'h8C51, 16'hA514, 16'hA554, 16'hA555, 16'h9492, 16'h934E, 16'h82CB, 16'hC555, 16'hDE59, 16'hACD3, 16'h5A48, 16'hA452, 16'hE65A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE1A, 16'hE61A, 16'hE65A, 16'hE61A, 16'hE619, 16'hE61A, 16'hDE19, 16'hDE19, 16'hD557, 16'hCD16, 16'hEE5B, 16'hDDD8, 16'hABD0, 16'h8A49, 16'hCC93, 16'hCCD4, 16'hCC93, 16'hCC94, 16'hBB8F, 16'hAB0D, 16'hDD16, 16'hE557, 16'hF5D9, 16'hF61A, 16'hF61A, 16'hF65B, 16'hFEDD, 16'hFEDD, 16'hFEDD, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF71D, 16'h6A09, 16'h5000, 16'h8187, 16'hCB0E, 16'hCB4F,
        16'hCB4F, 16'hCB0F, 16'hCB4F, 16'hCB0F, 16'hCB4F, 16'hE454, 16'hF4D6, 16'hECD5, 16'hEC95, 16'hEC95, 16'hEC95, 16'hECD5, 16'hEC95, 16'hEC95, 16'hECD5, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC54, 16'hE412, 16'hB1CA, 16'hCD56, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5F, 16'hEE9C, 16'h930D, 16'hE619, 16'hE65A, 16'hE65A, 16'hE619, 16'hEE5B, 16'hC4D4, 16'h8187, 16'h928B, 16'hDDD8, 16'hE65A, 16'hD5D8, 16'hD5D8, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD9, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD9, 16'hDE19, 16'hD597, 16'hCD56, 16'hD5D8, 16'hC515, 16'h51C7, 16'h8450, 16'h5A89, 16'hACD4, 16'hBD55, 16'hB515, 16'hB514, 16'hB514, 16'h8B4E, 16'hBD56, 16'hD618, 16'h6A4A, 16'h8C91, 16'hAD95, 16'h9D13, 16'h738E, 16'h94D2, 16'hAD95, 16'hA554, 16'h744F, 16'h6C0E, 16'h9D54, 16'hA595, 16'hA554, 16'hA595, 16'hA595, 16'hA555, 16'hA555,
        16'hA594, 16'h8450, 16'hAD55, 16'hAD95, 16'hC6DA, 16'hBE58, 16'hEF5D, 16'hFFDF, 16'hBD55, 16'h9C91, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h6289, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h6B4C, 16'h9D94, 16'h73CE, 16'hA4D2, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB555, 16'hD659, 16'hFFDF, 16'hBD56, 16'hA4D3, 16'hDE9A, 16'hCE58, 16'h730C, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h9C10, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE18, 16'h7B0C, 16'hCDD7, 16'hD619, 16'hD618, 16'hD618, 16'hD618, 16'hD659, 16'hB4D4, 16'hBD55, 16'hBD55, 16'h638D, 16'h9D54, 16'h9513, 16'h8CD2, 16'h8CD2, 16'h8491, 16'h8C91, 16'h9D13, 16'hAD54, 16'hA554, 16'hA554, 16'hA554, 16'h94D2, 16'h7C0F, 16'hA554, 16'hA554, 16'hA554, 16'h94D2, 16'h8B4E, 16'h830C, 16'hC555, 16'hDE59, 16'hAC93, 16'h5A48, 16'h9C10,
        16'hDE5A, 16'hDE1A, 16'hDE1A, 16'hDE19, 16'hE65A, 16'hE61A, 16'hE61A, 16'hE619, 16'hE619, 16'hE61A, 16'hDE19, 16'hDE19, 16'hD598, 16'hC4D5, 16'hE65A, 16'hE619, 16'h828A, 16'hAB4E, 16'hD515, 16'hCCD4, 16'hD4D4, 16'hCCD4, 16'hCC52, 16'hAACC, 16'hED98, 16'hEDD9, 16'hED98, 16'hED98, 16'hF598, 16'hF5D9, 16'hF61A, 16'hF69B, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hEEDC, 16'h5002, 16'h5800, 16'h9A0A, 16'hCB4F, 16'hCB4F, 16'hCB4F, 16'hCB4F, 16'hCB4F, 16'hCB0F, 16'hE454, 16'hF4D6, 16'hEC95, 16'hECD5, 16'hECD5, 16'hEC95, 16'hECD5, 16'hECD5, 16'hECD5, 16'hECD5, 16'hECD6, 16'hF4D6, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hF495, 16'hCACD, 16'hCD15, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF9F,
        16'hC515, 16'hB452, 16'hEE5B, 16'hE61A, 16'hE61A, 16'hE65A, 16'hDD98, 16'h92CB, 16'hB34E, 16'h934E, 16'hE61A, 16'hE65A, 16'hD5D8, 16'hD5D8, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD9, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD5D8, 16'hCD56, 16'hD597, 16'hD5D8, 16'h8B8E, 16'h6B8D, 16'h8450, 16'h6A8B, 16'hBD55, 16'hB515, 16'hB555, 16'hBD55, 16'hAC93, 16'h8B4D, 16'hD5D8, 16'hC555, 16'h5A08, 16'h9D13, 16'h8C91, 16'h7C50, 16'h9D54, 16'hA595, 16'hA555, 16'h9D54, 16'h6C0F, 16'h744F, 16'hA595, 16'hA555, 16'hA595, 16'hA595, 16'hA595, 16'hA595, 16'hA595, 16'h9513, 16'h8C51, 16'hBDD6, 16'hAD95, 16'hBED9, 16'hCE99, 16'hFFDF, 16'hFFDF, 16'hA492, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hB555, 16'h8C0F, 16'hFFDE, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h7BCE, 16'h8490, 16'h6B8D, 16'h9410, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hEF1C, 16'hACD3, 16'hF79E, 16'hFFDF, 16'hBD96, 16'h9C92, 16'hDE9A, 16'hAD14, 16'h838E, 16'hF79D, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h8BCF, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA492, 16'h93D0, 16'hD619, 16'hD618, 16'hCE18, 16'hCE18, 16'hCE18, 16'hD619, 16'h9C11, 16'hE65A, 16'h9C51, 16'h6BCE, 16'hA554, 16'h9D53, 16'h8CD2, 16'h8CD2, 16'h8CD1, 16'h8C91, 16'h9D13, 16'hAD54, 16'hA554, 16'hA554, 16'hAD95, 16'h8450, 16'h8450, 16'hAD95, 16'hA554, 16'hA554, 16'h94D2, 16'h8B4D, 16'h8B0C, 16'hBD14, 16'hDE5A, 16'hACD3, 16'h6ACA, 16'h8B8E, 16'hDE19, 16'hDE1A, 16'hDE1A, 16'hE65A, 16'hDE1A, 16'hE65A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hDE19, 16'hDE19, 16'hDDD8, 16'hC4D4, 16'hDDD9, 16'hEE5B, 16'h7ACB, 16'h92CC, 16'hD4D5, 16'hD515, 16'hD4D5, 16'hD4D4, 16'hD4D5, 16'hAACC, 16'hE556, 16'hFF1D, 16'hFF1D, 16'hFEDD, 16'hFEDD, 16'hFF1D, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hE69B, 16'h4800, 16'h6082, 16'hB28C, 16'hCB4F, 16'hCB0F, 16'hCB4F, 16'hCB4F, 16'hCB0F, 16'hE453, 16'hF4D6, 16'hEC95, 16'hECD5, 16'hEC95, 16'hECD5, 16'hECD6, 16'hECD5, 16'hECD6, 16'hECD6, 16'hECD6, 16'hF4D6, 16'hF4D6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hE391, 16'hDD56, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF1D, 16'h9B4E, 16'hDDD8, 16'hE65A, 16'hE61A, 16'hE65A, 16'hEE1A, 16'h930D, 16'hC411, 16'hA2CC, 16'hAC52, 16'hEE5A, 16'hDE19, 16'hD5D8, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD8, 16'hC556, 16'hCD97, 16'hD5D8, 16'hC515, 16'h49C7, 16'h9513, 16'h6B4C, 16'h93D0, 16'hBD56, 16'hBD55, 16'hBD55, 16'hBD56, 16'h9C10, 16'h9C10, 16'hDE19, 16'hAC92, 16'h630B, 16'h8C91, 16'h8C92, 16'hA595, 16'hA595,
        16'h9D54, 16'hA595, 16'h9D54, 16'h63CE, 16'h8491, 16'hA595, 16'hA595, 16'hA595, 16'hA595, 16'hA595, 16'hA595, 16'hADD6, 16'h8C91, 16'hA513, 16'hBD95, 16'hB5D6, 16'hB698, 16'hD6DB, 16'hFFDF, 16'hF75D, 16'h8BCE, 16'hE6DB, 16'hFFDF, 16'hEF5D, 16'h838C, 16'hDEDA, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD618, 16'h6ACA, 16'h4A89, 16'h4A89, 16'h9C91, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCDD7, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hC5D7, 16'h9C92, 16'hD659, 16'h8BCF, 16'hAD13, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79D, 16'h8B8E, 16'hDEDA, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79D, 16'h834D, 16'hB514, 16'hD619, 16'hCE18, 16'hD618, 16'hCE18, 16'hD659, 16'hBD56, 16'hA492, 16'hEEDC, 16'h7B4D, 16'h7C10, 16'hA594, 16'h9D54, 16'h8CD2, 16'h8CD2, 16'h8491, 16'h8CD2, 16'hA554, 16'hAD95, 16'hA554, 16'hA595, 16'hAD95, 16'h634D,
        16'h8450, 16'hAD95, 16'h9D54, 16'h9D54, 16'h9D13, 16'h834D, 16'h82CB, 16'hAC92, 16'hDE5A, 16'hB514, 16'h6B0B, 16'h7B4D, 16'hD5D8, 16'hDE5A, 16'hDE1A, 16'hDE1A, 16'hDE1A, 16'hDE19, 16'hE65A, 16'hE61A, 16'hE61A, 16'hE61A, 16'hDE19, 16'hDE19, 16'hE5D9, 16'hCCD5, 16'hD598, 16'hEE5B, 16'h8B8E, 16'h000, 16'h824A, 16'hB411, 16'hD4D5, 16'hDD15, 16'hDD56, 16'hBB90, 16'hBC11, 16'hFEDD, 16'hF71D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hEEDC, 16'h5000, 16'h7104, 16'hC30E, 16'hCB4F, 16'hCB4F, 16'hCB4F, 16'hCB0F, 16'hDBD2, 16'hF4D6, 16'hEC95, 16'hECD5, 16'hECD5, 16'hEC95, 16'hECD5, 16'hECD5, 16'hECD6, 16'hECD5, 16'hECD6, 16'hECD6, 16'hECD5, 16'hECD5, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD5, 16'hECD5, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC13, 16'hEDD9, 16'hFF9F,
        16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hD5D8, 16'hA38F, 16'hEE5B, 16'hE61A, 16'hE65A, 16'hEE5A, 16'hA38F, 16'hAB4E, 16'hDC94, 16'h8A09, 16'hCD97, 16'hE65A, 16'hD5D8, 16'hD5D8, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD9, 16'hDDD9, 16'hDDD9, 16'hDE19, 16'hDE19, 16'hDDD9, 16'hCD56, 16'hC556, 16'hD597, 16'hD5D8, 16'h830C, 16'h740F, 16'h9D54, 16'h5207, 16'hB514, 16'hBD56, 16'hBD55, 16'hBD56, 16'hBD55, 16'h7B0C, 16'hB514, 16'hD5D8, 16'h728B, 16'h8C91, 16'hADD6, 16'hA595, 16'hA595, 16'hA595, 16'hA595, 16'hA595, 16'h9513, 16'h63CE, 16'h9513, 16'hAD95, 16'hA595, 16'hA595, 16'hA595, 16'hA595, 16'hA595, 16'hA596, 16'h7C0F, 16'hBD96, 16'hB514, 16'hBE18, 16'hB617, 16'hEF5D, 16'hFFDF, 16'hD659, 16'h940F, 16'hFF9E, 16'hFFDF, 16'hACD3, 16'hB555, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hCE18, 16'h8BCF, 16'h000, 16'h3000, 16'h7B8D, 16'hC5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hB514, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h9451, 16'hC5D7, 16'h730B, 16'hD658, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h8B8E, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h7ACB, 16'hC597, 16'hD619, 16'hCE18, 16'hD618, 16'hCE18, 16'hD619, 16'h9C51, 16'hCDD8, 16'hE6DB, 16'h730C, 16'h8450, 16'hA595, 16'hA594, 16'h8CD2, 16'h8CD2, 16'h84D1, 16'h94D2, 16'hA554, 16'hA595, 16'hA555, 16'hAD95, 16'h9513, 16'h4248, 16'h8CD2, 16'hAD95, 16'h9D54, 16'h9D54, 16'h9D14, 16'h834D, 16'h830C, 16'hAC52, 16'hDE5A, 16'hB515, 16'h6B0B, 16'h730C, 16'hCD97, 16'hE65A, 16'hDE1A, 16'hDE1A, 16'hDE19, 16'hE65A, 16'hE65A, 16'hE61A, 16'hE61A, 16'hDE19, 16'hDE1A, 16'hDE19, 16'hE619, 16'hCCD5, 16'hD597, 16'hEE5B, 16'h8B8E, 16'h5289, 16'h528A, 16'h3041, 16'h7209, 16'hAB8F, 16'hCCD4, 16'hD453, 16'hA2CC, 16'hFE9B, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E,
        16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF71D, 16'h6186, 16'h8146, 16'hCB4F, 16'hCB0F, 16'hCB4F, 16'hCB0F, 16'hD390, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hF4D6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD5, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD5, 16'hECD5, 16'hECD6, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC54, 16'hF65B, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hA38F, 16'hD556, 16'hEE5A, 16'hE65A, 16'hEE5A, 16'hA3D0, 16'h9ACC, 16'hDD15, 16'hC412, 16'h82CB, 16'hE619, 16'hDE19, 16'hD5D9, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD9, 16'hDE19, 16'hDE19, 16'hCD57, 16'hC556, 16'hD597, 16'hDDD8, 16'hB493, 16'h49C6, 16'hA595, 16'h7C0F, 16'h72CB, 16'hC596, 16'hBD56,
        16'hBD55, 16'hBD56, 16'hAC93, 16'h728A, 16'hCDD8, 16'hC556, 16'h628A, 16'hA595, 16'hA595, 16'hA595, 16'hA595, 16'hA555, 16'hA595, 16'hAD95, 16'h8CD2, 16'h6C0E, 16'hA595, 16'hA595, 16'hA595, 16'hADD6, 16'hA595, 16'hA595, 16'hA595, 16'hA595, 16'h7C0F, 16'hC5D7, 16'hB555, 16'hB617, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hA4D2, 16'hC5D6, 16'hFFDF, 16'hD618, 16'hAD13, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD699, 16'hACD3, 16'hACD3, 16'hC5D6, 16'hDE9A, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hB514, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8C10, 16'hACD4, 16'h7B0B, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h8BCF, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC5D7, 16'h830C, 16'hD618, 16'hD619, 16'hCE18, 16'hCE18, 16'hD618, 16'hCDD8, 16'h8B8E, 16'hEF1C, 16'hCE58, 16'h9450, 16'h8450,
        16'hADD6, 16'hA595, 16'h8CD2, 16'h8CD2, 16'h8CD2, 16'h94D2, 16'hA554, 16'hA595, 16'hA595, 16'hAD95, 16'h8451, 16'h734D, 16'h94D2, 16'hADD5, 16'hA554, 16'h9D54, 16'hA554, 16'h838D, 16'h8B0C, 16'h9C10, 16'hDE19, 16'hBD96, 16'h6B0B, 16'h6B0B, 16'hBD14, 16'hE65A, 16'hDE19, 16'hDE1A, 16'hDE1A, 16'hDE1A, 16'hE65A, 16'hDE1A, 16'hDE19, 16'hDE1A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hCD16, 16'hCD56, 16'hEE5B, 16'h9C11, 16'h4A89, 16'h740F, 16'h6B8C, 16'h5A89, 16'h4185, 16'h5945, 16'h71C8, 16'h5800, 16'hDD97, 16'hFF1E, 16'hFF1D, 16'hFF1E, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'h7ACC, 16'h8146, 16'hD34F, 16'hCB0F, 16'hCB4F, 16'hCB4F, 16'hE453, 16'hF4D6, 16'hEC95, 16'hECD5, 16'hECD5, 16'hEC95, 16'hECD6, 16'hECD6, 16'hF4D6, 16'hECD6, 16'hF4D6, 16'hF4D6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hF4D6, 16'hF4D6, 16'hECD6, 16'hECD5,
        16'hECD6, 16'hECD6, 16'hECD6, 16'hECD5, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hEC95, 16'hE495, 16'hFF1D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hD597, 16'hA38F, 16'hEE1A, 16'hEE5B, 16'hE5D9, 16'h9B4E, 16'h9ACC, 16'hDCD5, 16'hE516, 16'hA30D, 16'h9BD0, 16'hEE5A, 16'hD5D9, 16'hDDD9, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hCD97, 16'hC556, 16'hCD97, 16'hD5D8, 16'hD5D8, 16'h6A89, 16'h8491, 16'hA595, 16'h4A08, 16'h9C51, 16'hC597, 16'hBD55, 16'hBD96, 16'hC597, 16'h830C, 16'h9410, 16'hDE19, 16'h93D0, 16'h73CE, 16'hADD6, 16'hA595, 16'hA595, 16'hA595, 16'hA595, 16'hA595, 16'hA595, 16'h7C91, 16'h7C50, 16'hADD6, 16'hA595, 16'hAD95, 16'hADD6, 16'hA595, 16'hA595, 16'hADD6, 16'h94D3, 16'h9491, 16'hC5D7, 16'hAD55, 16'hA554, 16'hEF5C, 16'hFFDF, 16'hE71B, 16'h838D, 16'hF75D, 16'hEF5D, 16'hC5D7, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'hC596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h8C10, 16'h8BCF, 16'h8BCE, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDE, 16'h8C0F, 16'hD618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hACD3, 16'h8BCF, 16'hD618, 16'hCE18, 16'hCE18, 16'hCE18, 16'hCE19, 16'hB514, 16'hA451, 16'hFF9E, 16'hC5D6, 16'hB554, 16'h7C50, 16'hADD6, 16'hA595, 16'h8D12, 16'h8CD2, 16'h84D2, 16'h94D2, 16'hA595, 16'hA595, 16'hAD96, 16'h9D14, 16'h9C92, 16'hA492, 16'h8CD1, 16'hADD5, 16'hA595, 16'hA554, 16'hA595, 16'h83CF, 16'h8B0D, 16'h8B8E, 16'hD5D8, 16'hCDD7, 16'h734C, 16'h6B0B, 16'hA452, 16'hDE19, 16'hDE19, 16'hDE59, 16'hDE1A, 16'hDE19, 16'hDE1A, 16'hDE1A, 16'hDE19, 16'hDE1A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD557, 16'hCD56, 16'hEE9B, 16'hAC92, 16'h4A89, 16'h740F, 16'h6BCD,
        16'h740E, 16'h73CD, 16'h6B8C, 16'h634C, 16'h4184, 16'hB3D0, 16'hFEDD, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'h9C11, 16'h8905, 16'hD350, 16'hCB4F, 16'hCB0E, 16'hD390, 16'hEC95, 16'hEC95, 16'hEC95, 16'hECD5, 16'hECD5, 16'hECD5, 16'hECD6, 16'hECD6, 16'hECD6, 16'hF4D6, 16'hECD6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hECD6, 16'hECD6, 16'hF4D6, 16'hECD5, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hF4D6, 16'hEC95, 16'hEC95, 16'hEC95, 16'hECD5, 16'hEC95, 16'hED17, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hF6DC, 16'h92CB, 16'hDDD8, 16'hF65B, 16'hDD57, 16'h8A8B, 16'hA34E, 16'hDCD5, 16'hE4D6, 16'hD493, 16'h4000, 16'hBCD4, 16'hE65A, 16'hDDD9, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD5D8,
        16'hCD97, 16'hD598, 16'hD5D8, 16'hE61A, 16'h9C11, 16'h52C9, 16'hA5D6, 16'h8C91, 16'h5A07, 16'hBD55, 16'hC596, 16'hBD56, 16'hC597, 16'hB4D3, 16'h6208, 16'hC596, 16'hCDD8, 16'h6A8A, 16'h9D14, 16'hA5D6, 16'hA595, 16'hA595, 16'hA596, 16'hA595, 16'hA595, 16'hA595, 16'h73CE, 16'h8491, 16'hADD6, 16'hAD95, 16'hAD95, 16'hAD96, 16'hAD95, 16'hA5D5, 16'hADD6, 16'h7C10, 16'hBD96, 16'hBD95, 16'h83CE, 16'hCE58, 16'hFFDF, 16'hFFDF, 16'hAD13, 16'hAD14, 16'hFFDF, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE18, 16'hCDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9451, 16'h6A8A, 16'hA492, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9C91, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9410,
        16'hA492, 16'hD659, 16'hCE18, 16'hCE18, 16'hCE18, 16'hCE18, 16'h9C10, 16'hC596, 16'hFF9E, 16'hBD95, 16'hCE18, 16'h7C0F, 16'hADD6, 16'hA595, 16'h9513, 16'h84D1, 16'h84D2, 16'h9513, 16'hA595, 16'hA595, 16'hADD6, 16'h7C50, 16'hBD96, 16'hB555, 16'h8491, 16'hAD95, 16'hA555, 16'hA555, 16'hA595, 16'h8C50, 16'h830C, 16'h834D, 16'hCDD7, 16'hD618, 16'h7B8D, 16'h6B4C, 16'h8B8F, 16'hDE19, 16'hDE59, 16'hDE59, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE1A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD598, 16'hCD97, 16'hE65A, 16'hBCD4, 16'h4A89, 16'h7C50, 16'h63CD, 16'h6BCD, 16'h6BCD, 16'h6BCD, 16'h740E, 16'h6B8D, 16'h6945, 16'hEE5A, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hCDD8, 16'h7800, 16'hD390, 16'hCB4F, 16'hCB4F, 16'hE453, 16'hECD5, 16'hEC95, 16'hEC95, 16'hEC95, 16'hECD5, 16'hF4D6, 16'hF4D6,
        16'hECD6, 16'hECD6, 16'hF4D6, 16'hECD6, 16'hECD6, 16'hF4D6, 16'hF4D6, 16'hECD6, 16'hF4D6, 16'hF4D6, 16'hECD6, 16'hF4D6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD5, 16'hECD5, 16'hECD5, 16'hECD6, 16'hEC54, 16'hEE19, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF5F, 16'hBC11, 16'hD4D5, 16'hEE1A, 16'hB411, 16'h8A4A, 16'hC411, 16'hE557, 16'hE557, 16'hE516, 16'h92CB, 16'h5186, 16'hD598, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD9, 16'hDE19, 16'hD5D8, 16'hCD97, 16'hD5D8, 16'hD5D8, 16'hDE19, 16'hC515, 16'h4186, 16'h9513, 16'hA5D6, 16'h630B, 16'h8BCF, 16'hC5D7, 16'hC597, 16'hC597, 16'hCDD7, 16'h7ACB, 16'h8BCF, 16'hDE59, 16'h93D0, 16'h73CE, 16'hADD6, 16'hA595, 16'hA5D6, 16'hA596, 16'hA596, 16'hA595, 16'hADD6, 16'h9D13, 16'h5B0B, 16'h8CD2, 16'hADD6, 16'hADD6, 16'hADD6, 16'hADD6, 16'hADD6, 16'hADD6, 16'hA595, 16'h8C0F, 16'hCDD7, 16'h838E, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hEF5C, 16'h7B4C, 16'hEF1C,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC5D7, 16'hD619, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD14, 16'h4080, 16'hB514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB555, 16'hA4D3, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h834D, 16'hACD4, 16'hD659, 16'hCE18, 16'hCE18, 16'hCE18, 16'hCDD8, 16'h834E, 16'hE6DB, 16'hF75E, 16'hBD96, 16'hDE9A, 16'h740F, 16'hADD6, 16'hA5D6, 16'h9513, 16'h84D2, 16'h84D1, 16'h9553, 16'hA595, 16'hA595, 16'hA596, 16'h6B8D, 16'hE6DB, 16'hB555, 16'h8491, 16'hADD6, 16'hA595, 16'hA595, 16'hA595, 16'h94D2, 16'h7ACB, 16'h7ACB, 16'hC597, 16'hD619, 16'h83CF, 16'h6B4C, 16'h7B8D, 16'hD5D8, 16'hDE59, 16'hDE19, 16'hDE1A, 16'hDE1A, 16'hDE1A, 16'hDE1A,
        16'hDE19, 16'hDE1A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD9, 16'hD597, 16'hDE1A, 16'hCD56, 16'h4A47, 16'h7C50, 16'h6C0E, 16'h6BCD, 16'h6BCD, 16'h6BCD, 16'h6BCD, 16'h740E, 16'h3984, 16'hBC92, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF71D, 16'h71C7, 16'hC30E, 16'hCB4F, 16'hD390, 16'hEC95, 16'hECD5, 16'hECD5, 16'hECD5, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hF4D6, 16'hECD6, 16'hF4D6, 16'hECD6, 16'hECD6, 16'hF4D6, 16'hF4D6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD5, 16'hECD6, 16'hECD6, 16'hF4D6, 16'hE413, 16'hF71D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hF71D, 16'hFF9F, 16'hFF5F, 16'hF6DC, 16'hB451, 16'hA2CC, 16'hBC12, 16'h92CC, 16'hB38F, 16'hDD16, 16'hEDD9, 16'hF5DA, 16'hF599, 16'hC412, 16'h5104, 16'h8B4E,
        16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hDE19, 16'hD597, 16'h61C8, 16'h7C50, 16'hA5D6, 16'h9513, 16'h5208, 16'hBD55, 16'hCDD7, 16'hC597, 16'hCDD8, 16'hAC92, 16'h61C7, 16'hC597, 16'hC556, 16'h51C7, 16'h9D54, 16'hADD6, 16'hA595, 16'hA596, 16'hA596, 16'hA595, 16'hA595, 16'hADD6, 16'h8C90, 16'h73CD, 16'h9513, 16'hAE16, 16'hADD6, 16'hADD6, 16'hADD6, 16'hADD6, 16'hADD6, 16'h94D2, 16'h8C0F, 16'hA491, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD13, 16'hB514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC596, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h2000,
        16'hBD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h838E, 16'hF79E, 16'hFFDF, 16'hEF5D, 16'h72CB, 16'hB555, 16'hD659, 16'hCE18, 16'hCE18, 16'hCE18, 16'hBD56, 16'h8B8E, 16'hF79E, 16'hEF1C, 16'hC5D7, 16'hE6DB, 16'h73CE, 16'hADD6, 16'hA5D6, 16'h9513, 16'h84D2, 16'h84D1, 16'h9D54, 16'hA595, 16'hADD6, 16'h9D54, 16'h83CE, 16'hFF9E, 16'hB555, 16'h8450, 16'hADD6, 16'hA595, 16'hA595, 16'hA595, 16'hA594, 16'h7B4C, 16'h728A, 16'hACD4, 16'hDE59, 16'h9C92, 16'h634B, 16'h6B4C, 16'hBD15, 16'hDE5A, 16'hDE19, 16'hDE19, 16'hDE1A, 16'hDE1A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD9, 16'hD5D8, 16'hDE19, 16'hDDD8, 16'h6A8A, 16'h740F, 16'h8491, 16'h73CE, 16'h6BCD, 16'h6BCE, 16'h740E, 16'h740F, 16'h6B8D, 16'h6987, 16'hF69B, 16'hFF1E, 16'hFF1D, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF,
        16'hB4D4, 16'h9947, 16'hD390, 16'hD3D1, 16'hECD5, 16'hECD5, 16'hEC95, 16'hEC95, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hF4D6, 16'hF4D6, 16'hECD6, 16'hECD6, 16'hF4D6, 16'hF4D6, 16'hECD6, 16'hECD6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hECD6, 16'hF4D6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hF4D6, 16'hECD5, 16'hF4D6, 16'hEC54, 16'hE5D9, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hDDD9, 16'hC4D3, 16'hBC11, 16'h9A8A, 16'h9249, 16'hB3D0, 16'hC452, 16'hE557, 16'hEDD9, 16'hF65C, 16'hFE9D, 16'hFE5C, 16'hD4D4, 16'h5985, 16'h59C7, 16'hACD3, 16'hE65A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD9, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hDDD8, 16'hDE19, 16'h7B0C, 16'h5B4C, 16'h9D95, 16'hA5D6, 16'h634C, 16'h93CF, 16'hCDD7, 16'hC597, 16'hCDD7, 16'hBD15, 16'h5945, 16'hAC93, 16'hCDD7, 16'h6249, 16'h8450, 16'hADD6, 16'hA596, 16'hA596, 16'hA596, 16'hA596, 16'hAD96, 16'hADD6, 16'hA555, 16'h840F, 16'h9D12, 16'h9513, 16'hB617, 16'hADD6, 16'hADD6, 16'hADD6,
        16'hADD6, 16'hADD6, 16'h738D, 16'h9C92, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h838E, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD96, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h4080, 16'hBD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h7B4D, 16'hDEDB, 16'hFFDF, 16'hE71C, 16'h6A8A, 16'hBD96, 16'hD619, 16'hCE18, 16'hCE18, 16'hD659, 16'hACD3, 16'hAC93, 16'hFFDF, 16'hE69B, 16'hC5D7, 16'hEF5D, 16'h738D, 16'hA595, 16'hADD6, 16'h9554, 16'h84D2, 16'h84D2, 16'h9D54, 16'hA595, 16'hADD6, 16'h8C92, 16'hA4D2, 16'hFFDF, 16'hB555, 16'h7C50, 16'hADD6, 16'hA595, 16'hA595, 16'hA595, 16'hA595, 16'h83CE, 16'h7A8B,
        16'h9C51, 16'hDE59, 16'hBD96, 16'h5289, 16'h5ACA, 16'h9C51, 16'hDE5A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE1A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD5D8, 16'hDDD9, 16'hE61A, 16'h938F, 16'h638C, 16'h9554, 16'h8492, 16'h7C50, 16'h7C50, 16'h8491, 16'h8491, 16'h8CD1, 16'h4A88, 16'hB411, 16'hFEDE, 16'hFF1D, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF71D, 16'h8248, 16'hC30E, 16'hE412, 16'hECD5, 16'hEC95, 16'hEC95, 16'hF4D6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hEC95, 16'hE516, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF71D, 16'hEEDB, 16'hF6DB,
        16'hFEDC, 16'hFEDC, 16'hFF1D, 16'hFF1E, 16'hFF1E, 16'hFF1F, 16'hFEDE, 16'hDD16, 16'h5945, 16'h7B4C, 16'h728A, 16'hD5D8, 16'hE65A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD9, 16'hD5D8, 16'hD5D8, 16'hDE19, 16'h93CF, 16'h528A, 16'h9D54, 16'hA5D6, 16'h84D1, 16'h6249, 16'hC596, 16'hC5D7, 16'hCDD8, 16'hC556, 16'h6A08, 16'h9C11, 16'hCD97, 16'h728A, 16'h738E, 16'hADD6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hADD6, 16'hA595, 16'hADD6, 16'h8451, 16'hAD13, 16'hAD54, 16'h9D54, 16'hB617, 16'hADD6, 16'hADD6, 16'hADD6, 16'hADD7, 16'h9D54, 16'h6B0B, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h72CA, 16'hDE99, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCDD7, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h6A8A, 16'hBD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9C92, 16'hB554, 16'hFFDF, 16'hDE9A, 16'h6A49, 16'hC5D7, 16'hCE19, 16'hCE18, 16'hCE18, 16'hCE18, 16'h9C10, 16'hCDD8, 16'hFFDF, 16'hDE9A, 16'hC5D7, 16'hF79E, 16'h7BCE, 16'hA595, 16'hB617, 16'h9D94, 16'h84D2, 16'h8CD2, 16'h9D94, 16'hADD6, 16'hAE16, 16'h73CE, 16'hCDD7, 16'hFFDF, 16'hBDD6, 16'h7C0F, 16'hAE16, 16'hA5D5, 16'hA595, 16'hA595, 16'hAD96, 16'h9492, 16'h728B, 16'h8B8E, 16'hCDD8, 16'hD618, 16'h7B4D, 16'h5289, 16'h734C, 16'hD618, 16'hDE19, 16'hDE19, 16'hDE5A, 16'hDE5A, 16'hDE19, 16'hDE1A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD5D9, 16'hE61A, 16'hB4D4, 16'h5289, 16'h9D14, 16'h9514, 16'h8D13, 16'h8CD2, 16'h8CD2, 16'h84D1, 16'h84D1, 16'h7C4F, 16'h4040, 16'hDD57, 16'hFF1E, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hD618, 16'h8000, 16'hE412, 16'hF4D5, 16'hECD5, 16'hECD5, 16'hECD6, 16'hECD6, 16'hECD5, 16'hECD6, 16'hF4D6, 16'hECD6, 16'hECD6, 16'hF4D6, 16'hF516, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hECD6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hF4D6, 16'hF4D6, 16'hDC54, 16'hF71D, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF1E, 16'hCD15, 16'h5800, 16'h7BCE, 16'h6B4C, 16'h9BD0, 16'hE65A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD5D8, 16'hE65A, 16'hA451, 16'h41C6, 16'h9513, 16'h9DD5, 16'h9595, 16'h4A48, 16'hAC93, 16'hCDD7, 16'hCDD7, 16'hC556, 16'h6A8A, 16'h93D0, 16'hBD15, 16'h6248, 16'h6B4C, 16'hAD96, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hA5D6,
        16'hA5D6, 16'hA596, 16'hADD6, 16'hA5D6, 16'h5B0A, 16'hD699, 16'h9CD2, 16'h9D95, 16'hAE17, 16'hAE16, 16'hADD6, 16'hADD6, 16'hADD7, 16'h73CE, 16'hBD95, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DA, 16'h72C9, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9B, 16'hA493, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9C51, 16'hACD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h7B4C, 16'hFFDE, 16'hDE9A, 16'h6249, 16'hC5D7, 16'hCE18, 16'hCE18, 16'hCE18, 16'hCDD7, 16'h938E, 16'hE6DB, 16'hFFDF, 16'hDE9A, 16'hC597, 16'hFFDF, 16'h8C50, 16'h9513, 16'hB617, 16'hA595, 16'h84D1, 16'h84D2, 16'h9D95, 16'hB5D6, 16'hADD6,
        16'h6B4C, 16'hE71C, 16'hFFDF, 16'hCE18, 16'h7C0F, 16'hADD6, 16'hA595, 16'hA595, 16'hA595, 16'hA595, 16'hA554, 16'h7B4D, 16'h7ACB, 16'hBD15, 16'hDE5A, 16'hA492, 16'h5288, 16'h5A89, 16'hBD55, 16'hDE5A, 16'hDE19, 16'hDE5A, 16'hDE19, 16'hDE19, 16'hDE1A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD9, 16'hDDD9, 16'hDE19, 16'hD597, 16'h5A08, 16'h8C91, 16'h9D54, 16'h9513, 16'h9513, 16'h8D13, 16'h8CD2, 16'h8D12, 16'h8491, 16'h6BCE, 16'h6A49, 16'hF69B, 16'hFF1E, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hB493, 16'hA1C9, 16'hF4D6, 16'hECD5, 16'hECD6, 16'hECD6, 16'hECD6, 16'hF4D6, 16'hECD6, 16'hECD6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hECD6, 16'hF516, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hECD6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hE454, 16'hF69B, 16'hFFDF,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF5E, 16'hC4D4, 16'h3000, 16'h738C, 16'h8450, 16'h49C6, 16'hC556, 16'hDE5A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD9, 16'hDDD8, 16'hDE19, 16'hE65A, 16'hAC93, 16'h41C7, 16'h9553, 16'hA5D6, 16'hA5D5, 16'h5B8C, 16'h8B4E, 16'hCDD7, 16'hCDD7, 16'hB515, 16'h6209, 16'h8B8E, 16'hA452, 16'h59C6, 16'h7C0F, 16'hADD6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hADD6, 16'hADD6, 16'hADD6, 16'hAE17, 16'h7C0F, 16'h7BCE, 16'hEF1B, 16'h8410, 16'hA5D6, 16'hAE17, 16'hAE16, 16'hADD6, 16'hAE17, 16'h9D14, 16'h734C, 16'hF79D, 16'hFFDF, 16'hFF9E, 16'hC595, 16'h6A47, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hACD3, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC596, 16'hAC92, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h8BCF, 16'hCE18, 16'hD659, 16'h6248, 16'hCDD7, 16'hCE18, 16'hCE18, 16'hCE19, 16'hC597, 16'h8B4E, 16'hEF1C, 16'hFFDF, 16'hDE9A, 16'hC596, 16'hFFDF, 16'hA514, 16'h8450, 16'hB617, 16'hA5D5, 16'h84D2, 16'h8512, 16'hA595, 16'hADD6, 16'h9D54, 16'h7B8D, 16'hF79E, 16'hFFDF, 16'hD699, 16'h73CE, 16'hADD6, 16'hA596, 16'hA595, 16'hA595, 16'hA595, 16'hAD95, 16'h9491, 16'h5186, 16'h9C10, 16'hDE5A, 16'hC597, 16'h5A8A, 16'h4A07, 16'h8BCF, 16'hD618, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD5D8, 16'hDE19, 16'h938F, 16'h5B0B, 16'h9D54, 16'h9513, 16'h9513, 16'h8D13, 16'h8D13, 16'h9513, 16'h7C91, 16'h84D2,
        16'h73CF, 16'h8ACC, 16'hFEDC, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hBCD4, 16'hD34F, 16'hF4D6, 16'hECD6, 16'hECD6, 16'hECD6, 16'hF4D6, 16'hF4D6, 16'hECD6, 16'hECD6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF516, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hE454, 16'hEE5B, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF1E, 16'hB411, 16'h1800, 16'h62CA, 16'h844F, 16'h6B4C, 16'h728A, 16'hDE18, 16'hDE59, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE61A, 16'hB493, 16'h3984, 16'h8D13, 16'h9DD6, 16'hA5D6, 16'h740F, 16'h72CB, 16'hCD97, 16'hC556, 16'hA451,
        16'h5986, 16'h724A, 16'h7ACB, 16'h4A07, 16'h94D2, 16'hADD6, 16'hADD6, 16'hADD6, 16'hADD6, 16'hADD6, 16'hA5D6, 16'hADD6, 16'hADD6, 16'hAE17, 16'h9D13, 16'h800, 16'hBD96, 16'hE6DB, 16'h73CE, 16'hAE57, 16'hAE17, 16'hAE16, 16'hAE16, 16'hB617, 16'h6B8D, 16'hACD3, 16'hEF1C, 16'hC596, 16'h9C0F, 16'h93CE, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'hBD96, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h9C0F, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDA, 16'h8C0F, 16'h9410, 16'h6289, 16'hC5D7, 16'hCE18, 16'hCE18, 16'hCE19, 16'hBD55, 16'h93CF, 16'hFF9E, 16'hFFDF,
        16'hE69B, 16'hBD55, 16'hFFDF, 16'hC618, 16'h740E, 16'hB617, 16'hADD6, 16'h8512, 16'h8512, 16'hA595, 16'hB617, 16'h8C92, 16'h9450, 16'hFFDF, 16'hFFDF, 16'hDEDA, 16'h738D, 16'hADD6, 16'hADD6, 16'hA596, 16'hA595, 16'hA595, 16'hA595, 16'hA595, 16'h6B0C, 16'h6A8B, 16'hCDD7, 16'hDE5A, 16'h8BD0, 16'h4A47, 16'h628A, 16'hBD55, 16'hD619, 16'hDE19, 16'hDE59, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hCD97, 16'hDE19, 16'hC556, 16'h4986, 16'h8CD2, 16'h9513, 16'h8D13, 16'h8D13, 16'h8D13, 16'h9553, 16'h84D2, 16'h7C91, 16'h9D94, 16'h534C, 16'h934E, 16'hFEDC, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hE5D9, 16'hDC53, 16'hEC95, 16'hF4D6, 16'hECD6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hECD6,
        16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hEC95, 16'hE516, 16'hF69C, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hEE9B, 16'h8B0D, 16'h3984, 16'h5ACA, 16'h6B8D, 16'h8450, 16'h5185, 16'hB4D3, 16'hDE5A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE619, 16'hA451, 16'h4A07, 16'h8D53, 16'hA616, 16'hA5D5, 16'h740F, 16'h72CB, 16'hBD14, 16'hAC92, 16'h59C8, 16'h000, 16'h5248, 16'h6B4C, 16'h4247, 16'h9513, 16'hAE17, 16'hA5D6, 16'hADD6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hADD6, 16'hAE17, 16'h9D54, 16'h734D, 16'h6A49, 16'hEF1C, 16'hBD96, 16'h8450, 16'hB657, 16'hAE16, 16'hAE16, 16'hAE17, 16'h94D2, 16'h730B, 16'hEF1C, 16'hE6DB, 16'hD618, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'h940F, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h628A, 16'h5208, 16'hC596, 16'hCE18, 16'hCDD8, 16'hD659, 16'hB514, 16'h9C10, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hB514, 16'hFFDF, 16'hE71C, 16'h738D, 16'hA5D6, 16'hAE16, 16'h8D53, 16'h8D13, 16'hA5D5, 16'hB617, 16'h7BCF, 16'hAD14, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h738D, 16'hA5D6, 16'hADD6, 16'hA595, 16'hA595, 16'hA595, 16'hA595, 16'hA596, 16'h94D2, 16'h49C7, 16'hA4D3, 16'hDE5A, 16'hBD96, 16'h628A, 16'h3101, 16'hA492, 16'hCD97, 16'hD5D8, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19,
        16'hCD97, 16'hC556, 16'hE65A, 16'h8B4E, 16'h5B4C, 16'h9D54, 16'h9513, 16'h8D13, 16'h8D13, 16'h9554, 16'h8D12, 16'h7C91, 16'h8D54, 16'h9D94, 16'h738D, 16'h7A09, 16'hE61A, 16'hFF9F, 16'hFF9E, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hF71D, 16'hE516, 16'hEC94, 16'hF4D5, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF4D6, 16'hF516, 16'hF516, 16'hF516, 16'hF516, 16'hF516, 16'hF516, 16'hF516, 16'hF516, 16'hF4D6, 16'hF4D6, 16'hECD6, 16'hED16, 16'hEE1A, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hCD56, 16'h6144, 16'h630B, 16'h6B8D, 16'h4A89, 16'h8450, 16'h6B4C, 16'h728A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDDD8,
        16'h8B4E, 16'h5288, 16'h9D94, 16'hA5D6, 16'h8D13, 16'h5B0B, 16'h38C2, 16'h834D, 16'h6ACB, 16'h4A89, 16'h6C0E, 16'h8CD2, 16'h9D54, 16'h740E, 16'h638C, 16'hA5D6, 16'hADD6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hAE17, 16'h9513, 16'h8C0F, 16'hA451, 16'hACD3, 16'hFF9E, 16'h83CE, 16'h9D95, 16'hB657, 16'hAE17, 16'hAE17, 16'hADD6, 16'h5A88, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB514, 16'hBD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hD659, 16'h51C7, 16'hBD96, 16'hCE18, 16'hC5D7, 16'hCE59, 16'hA493, 16'hA492, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hB514, 16'hFF9E, 16'hFFDF, 16'h8C50, 16'h9513, 16'hB617, 16'h9554, 16'h8D12, 16'hA595, 16'hBE17, 16'h738E, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hF79D, 16'h7BCE, 16'h9D94, 16'hADD6, 16'hAD96, 16'hADD6, 16'hA595, 16'hA595, 16'hA596, 16'hAD96, 16'h73CE, 16'h5A49, 16'hCE18, 16'hDE59, 16'hA492, 16'h000, 16'h838E, 16'hC597, 16'hCD97, 16'hD619, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD619, 16'hAC93, 16'hDDD8, 16'hCD97, 16'h4146, 16'h8491, 16'h9D54, 16'h9554, 16'h8D13, 16'h9553, 16'h8D13, 16'h84D2, 16'h9554, 16'h9554, 16'h9D95, 16'h740F, 16'h6186, 16'hDDD8, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF65B,
        16'hED58, 16'hECD6, 16'hEC96, 16'hEC96, 16'hF4D6, 16'hF4D6, 16'hF517, 16'hF517, 16'hF4D6, 16'hF517, 16'hF516, 16'hF516, 16'hF516, 16'hF4D6, 16'hED17, 16'hED98, 16'hF65B, 16'hFF1E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hF6DC, 16'hA38F, 16'h3080, 16'h73CD, 16'h844F, 16'h5B0B, 16'h6B8C, 16'h840F, 16'h4986, 16'hBD14, 16'hE65A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE65A, 16'hC556, 16'h6A09, 16'h4A48, 16'h9D95, 16'h9554, 16'h6BCD, 16'h4247, 16'h4248, 16'h52CA, 16'h638D, 16'h8D12, 16'h9DD5, 16'hA5D6, 16'hA616, 16'h8CD2, 16'h634B, 16'h8491, 16'hAE16, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hADD6, 16'hADD6, 16'hA5D6, 16'hAE17, 16'h9513, 16'h83CF, 16'hE65A, 16'h93CF, 16'hE6DB, 16'hE6DB, 16'h73CD, 16'hB657, 16'hAE57, 16'hAE57, 16'hAE17, 16'h5ACA, 16'hB555, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h7ACB, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h6A8A, 16'hB555, 16'hCE18, 16'hC617, 16'hCE58, 16'h9C51, 16'hACD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB514, 16'hEF5D, 16'hFFDF, 16'hC618, 16'h6B8D, 16'hB617, 16'h9D95, 16'h8D13, 16'hA595, 16'hB617, 16'h630C, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9450, 16'h9512, 16'hAE17, 16'hA596, 16'hADD6, 16'hA5D5, 16'hA595, 16'hA596, 16'hA595, 16'hA595, 16'h630B, 16'h8C0F, 16'hDE5A, 16'hD5D8, 16'h6ACB, 16'h28C2,
        16'hB515, 16'hCDD7, 16'hCDD7, 16'hD619, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD619, 16'hD619, 16'hDE5A, 16'hAC92, 16'h8B8F, 16'hE65A, 16'hAC92, 16'h4207, 16'h9D54, 16'h9D54, 16'h9554, 16'h9554, 16'h9513, 16'h84D2, 16'h9554, 16'h9554, 16'h9554, 16'h9D95, 16'h8CD2, 16'h38C3, 16'h9BD0, 16'hF6DC, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF1E, 16'hF65B, 16'hF599, 16'hED58, 16'hED17, 16'hED16, 16'hED17, 16'hED17, 16'hED17, 16'hF517, 16'hF558, 16'hF5D9, 16'hF65B, 16'hFEDC, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF5E, 16'hD597, 16'h61C7, 16'h4206, 16'h7C0F, 16'h7C0F, 16'h73CD, 16'h5B0B, 16'h7C0F, 16'h5A89, 16'h8B4D,
        16'hDE59, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hAC92, 16'h5A08, 16'h6ACB, 16'h8490, 16'hA5D6, 16'h9D95, 16'h9513, 16'h9D94, 16'h9D94, 16'h7C90, 16'h9D95, 16'hA5D6, 16'hA5D5, 16'hA5D6, 16'h9553, 16'h7C0F, 16'h9C92, 16'h9553, 16'hAE17, 16'hA5D6, 16'hADD6, 16'hADD6, 16'hADD6, 16'hA5D6, 16'hAE17, 16'h9D13, 16'h6B0C, 16'hEEDB, 16'hC556, 16'h9C51, 16'hFFDF, 16'hA4D3, 16'h9513, 16'hB658, 16'hAE57, 16'hAE17, 16'h6B8C, 16'h9C91, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA452, 16'h93D0, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h730C, 16'hA4D3, 16'hCE18, 16'hC618, 16'hCE59, 16'h9C51, 16'hACD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC596, 16'hE6DA, 16'hFFDF, 16'hF75D, 16'h738D, 16'h9D54, 16'hAE16, 16'h8D13, 16'hA595, 16'hB617, 16'h5ACA, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD14, 16'h7C50, 16'hB617, 16'hADD6, 16'hA596, 16'hA5D5, 16'hA595, 16'hA5D6, 16'hA5D6, 16'hADD6, 16'hA555, 16'h4A48, 16'h9451, 16'hDE9A, 16'hC556, 16'h2000, 16'h83CE, 16'hCDD7, 16'hC5D7, 16'hCDD7, 16'hD619, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD619, 16'hD619, 16'hD619, 16'hDE19, 16'hBD15, 16'h000, 16'h93CF, 16'hDE19, 16'h834E, 16'h5B4C, 16'h9D55, 16'h9554, 16'h9554, 16'h9D54, 16'h84D2, 16'h8D13, 16'h9554, 16'h9554, 16'h9554, 16'h9554, 16'h9513, 16'h5ACA, 16'h7186, 16'hCD97, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hFEDD, 16'hF6DD, 16'hFEDD, 16'hFF1D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hEE9B, 16'hA3D0, 16'h1800, 16'h634C, 16'h7C4F, 16'h740E, 16'h7C0F, 16'h634C, 16'h6B8C, 16'h738D, 16'h6208, 16'hD5D7, 16'hDE5A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hD619, 16'hDE19, 16'hE619, 16'hCD96, 16'h8B8E, 16'h000, 16'hB554, 16'h9450, 16'h8D13, 16'hA5D6, 16'hA5D5, 16'hA5D6, 16'hA5D6, 16'h9594, 16'h7C91, 16'hA5D6, 16'h9DD5, 16'h9DD5, 16'hA5D5, 16'h73CE, 16'hC596, 16'hA492, 16'h9D94, 16'hAE17, 16'hA5D6, 16'hADD6, 16'hAE16, 16'hAE16, 16'hAE17, 16'h9513, 16'h5AC9, 16'hE69B, 16'hDE59, 16'h728A, 16'hF75D, 16'hF75D, 16'h83CE, 16'hAE16, 16'hAE57, 16'hAE16,
        16'h6B4C, 16'h83CE, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h728A, 16'hA451, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9410, 16'h9410, 16'hCE58, 16'hC618, 16'hCE58, 16'h9C51, 16'hACD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'hCDD7, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h638D, 16'hAE16, 16'h9554, 16'h9D95, 16'hB617, 16'h62CA, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h738D, 16'hAE16, 16'hADD6,
        16'hA5D6, 16'hA595, 16'hA595, 16'hA595, 16'hA5D6, 16'hA596, 16'hADD6, 16'h9513, 16'h39C6, 16'h9410, 16'hDE5A, 16'hACD3, 16'h000, 16'hB515, 16'hCE18, 16'hCDD7, 16'hCDD8, 16'hD619, 16'hD619, 16'hD619, 16'hD619, 16'hD619, 16'hDE19, 16'hD619, 16'hDE19, 16'hC556, 16'h6B4C, 16'h5ACB, 16'h7B4D, 16'hC555, 16'h628A, 16'h73CF, 16'h9D95, 16'h9554, 16'h9554, 16'h84D2, 16'h8D13, 16'h9594, 16'h9554, 16'h9554, 16'h9554, 16'h9D55, 16'hA595, 16'h73CF, 16'h3040, 16'h930D, 16'hDDD9, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF1D, 16'hCD15,
        16'h6881, 16'h3800, 16'h630A, 16'h7C4F, 16'h740E, 16'h740E, 16'h7C0E, 16'h634C, 16'h738D, 16'h3081, 16'hB514, 16'hE65A, 16'hDE19, 16'hDE19, 16'hDE19, 16'hDE19, 16'hE65A, 16'hD5D8, 16'hA411, 16'h6208, 16'h800, 16'h9C51, 16'hE69A, 16'h6B8D, 16'hA5D6, 16'h9DD5, 16'hA5D5, 16'h9DD5, 16'hA616, 16'h8491, 16'h744F, 16'hA5D6, 16'hA5D6, 16'hAE16, 16'h740F, 16'hB554, 16'hE69A, 16'h7BCE, 16'hADD6, 16'hA5D6, 16'hAE17, 16'hADD6, 16'hADD6, 16'hAE17, 16'h84D2, 16'h6ACA, 16'hEEDB, 16'hEE9B, 16'h830C, 16'hDE9A, 16'hFFDF, 16'hACD3, 16'h8491, 16'hBE98, 16'hA595, 16'h5ACA, 16'h8C0F, 16'hF79D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h8B8E, 16'h830C, 16'hCDD7, 16'hE6DB, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD55, 16'h6A8A, 16'hC5D7, 16'hC618, 16'hCE58, 16'hA492, 16'hA492, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hACD3, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h7B8D, 16'h84D2, 16'hA5D6, 16'h9D94, 16'hB617, 16'h62CA, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h7B8D, 16'hA595, 16'hADD7, 16'hADD6, 16'hA596, 16'h9D54, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'h9514, 16'h5289, 16'h7B8E, 16'hCD97, 16'h834D, 16'h730D, 16'hCE18, 16'hCDD8, 16'hCDD8, 16'hCDD8, 16'hD619, 16'hD659, 16'hD619, 16'hD619, 16'hD619, 16'hD619, 16'hDE19, 16'hD5D8, 16'h734D, 16'h9D54, 16'h740F, 16'h5A49, 16'h7ACC, 16'h2840, 16'h73CE, 16'h9514, 16'h9D95, 16'h9554, 16'h9553, 16'h9594, 16'h9554, 16'h9D54, 16'h9D54, 16'h9D54, 16'h9554, 16'h9D95,
        16'h9513, 16'h4A89, 16'h40C0, 16'h8B8E, 16'hDE19, 16'hFF5F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF5F, 16'hE5D9, 16'h928B, 16'h6000, 16'h9147, 16'h70C5, 16'h5B4B, 16'h7C4F, 16'h740E, 16'h740E, 16'h73CE, 16'h630B, 16'h28C2, 16'h9C51, 16'hDE59, 16'hDE59, 16'hDE19, 16'hDE19, 16'hDE1A, 16'hD5D8, 16'hAC52, 16'h6208, 16'h5A89, 16'h83CE, 16'h5A08, 16'hF75D, 16'hC596, 16'h740F, 16'hAE16, 16'h9DD5, 16'hA5D5, 16'hA5D6, 16'h9D94, 16'h4208, 16'h7C50, 16'hA5D6, 16'hAE16, 16'h8491, 16'h9450, 16'hFF9E, 16'hB555, 16'h8490, 16'hB657, 16'hAE17, 16'hAE16, 16'hAE17, 16'hAE17, 16'h7C50,
        16'h838D, 16'hEEDC, 16'hDE19, 16'h8B0C, 16'hD659, 16'hFFDF, 16'hDE9A, 16'h73CE, 16'hAE17, 16'h8CD2, 16'h5208, 16'hAD13, 16'hFFDE, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hD659, 16'hBD96, 16'hCE18, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h51C6, 16'hAD14, 16'hCE18, 16'hCE58, 16'hA4D3, 16'h9C51, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB514, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h4A48,
        16'h8491, 16'hA595, 16'hB617, 16'h6B4C, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h8C10, 16'h9513, 16'hAE17, 16'hADD6, 16'hA5D6, 16'h8CD2, 16'hA595, 16'hADD7, 16'hA5D6, 16'hADD6, 16'hA5D6, 16'hADD6, 16'hA5D6, 16'h73CE, 16'h5A89, 16'h938E, 16'h5186, 16'h9C52, 16'hD618, 16'hCDD8, 16'hCDD8, 16'hD618, 16'hD619, 16'hD619, 16'hD619, 16'hD619, 16'hD619, 16'hD619, 16'hDE19, 16'h8BCF, 16'h8451, 16'hAE17, 16'h9513, 16'h638D, 16'h4A48, 16'h000, 16'h1881, 16'h5B0B, 16'h740F, 16'h84D1, 16'h9554, 16'h9594, 16'h9554, 16'h9D54, 16'h9554, 16'h9554, 16'h9554, 16'h9D95, 16'h8CD2, 16'h8491, 16'h6B8D, 16'h4943, 16'h8B4D, 16'hD5D7, 16'hF71D, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF6DC, 16'hB410, 16'h6800, 16'h8843, 16'hB24A, 16'hC30D, 16'h7105, 16'h5B0B, 16'h7C0F, 16'h7C0F, 16'h7C4F, 16'h5ACA, 16'h000, 16'h9C10, 16'hDE59, 16'hE69A, 16'hE69A, 16'hDE19, 16'hC556, 16'h9C10, 16'h6248, 16'h5A89, 16'h8C92, 16'hA554, 16'h4185, 16'hCE18, 16'hFFDF, 16'h838D, 16'h9553, 16'hA5D6, 16'h9D95, 16'hA616, 16'h9D95, 16'h7B8D, 16'h730C, 16'h8CD2, 16'hAE17, 16'h8492, 16'h83CE, 16'hF79E, 16'hF75D, 16'h7B8E, 16'h9D95, 16'hAE17, 16'hAE17, 16'hAE57, 16'hAE17, 16'h6B8E, 16'h9450, 16'hE69A, 16'hC596, 16'hA451, 16'hEEDB, 16'hFFDF, 16'hF75D, 16'h7B8D, 16'h6BCE, 16'h6B8D, 16'h940F, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h8BCF, 16'h7B4D, 16'hCE18, 16'hCE58, 16'hAD13, 16'h8BCF, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hA492, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hD699, 16'h62CB, 16'h634B, 16'h8CD2, 16'h630B, 16'hC5D6, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB555, 16'h740F, 16'hAE17, 16'hAE17, 16'hAE17, 16'h7C50, 16'h8CD2, 16'hAE17, 16'hA5D6, 16'hA5D6, 16'hADD6, 16'hA5D6, 16'hA616, 16'hADD6, 16'h9514, 16'h73CE, 16'h5248, 16'h000, 16'hB514, 16'hD619, 16'hCDD8, 16'hCE18, 16'hD618, 16'hD618, 16'hD618, 16'hD619, 16'hD619, 16'hD619, 16'hDE19, 16'hAC93, 16'h630B, 16'hA5D5, 16'h9D96, 16'h9D95, 16'h9553,
        16'h84D2, 16'h7C50, 16'h7410, 16'h8491, 16'h84D2, 16'h9D95, 16'h9D94, 16'h9D54, 16'h9554, 16'h9D54, 16'h9D54, 16'h9554, 16'h9D54, 16'h9513, 16'h8492, 16'h9D55, 16'h9D54, 16'h740F, 16'h3142, 16'h61C7, 16'hA451, 16'hD5D8, 16'hF71D, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFEDD, 16'hCD15, 16'h8905, 16'h8000, 16'hB20A, 16'hC2CD, 16'hD3D0, 16'hD452, 16'h7186, 16'h6B8C, 16'h7C10, 16'h73CE, 16'h4247, 16'h4986, 16'hB514, 16'hE69A, 16'hDE5A, 16'hCD97, 16'hA451, 16'h72CB, 16'h5A08, 16'h634C, 16'h9512, 16'hADD6, 16'hA555, 16'h41C6, 16'hAD95, 16'hFFDF, 16'hD659, 16'h6B4B, 16'hA5D6, 16'hA5D5, 16'hA616, 16'h9D95, 16'h638C, 16'hD618, 16'hB514, 16'h9D95, 16'h8CD2,
        16'h838D, 16'hF75D, 16'hFFDF, 16'hC5D6, 16'h7C4F, 16'hAE57, 16'hAE17, 16'hAE57, 16'hA5D6, 16'h5B0B, 16'hAD13, 16'hFFDE, 16'hF79E, 16'hE6DB, 16'hFF9E, 16'hFF9E, 16'hD659, 16'h730B, 16'h5A89, 16'hA492, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h3000, 16'hACD3, 16'hCE58,
        16'hBD95, 16'h7B0C, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'hB514, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hBD95, 16'h9C91, 16'h628A, 16'hAD13, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDA, 16'h634C, 16'hADD7, 16'hAE17, 16'hAE17, 16'h7C50, 16'h6B8D, 16'hA5D6, 16'hA5D6, 16'hADD6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hAE17, 16'hADD7, 16'hA595, 16'h7C0F, 16'h4A07, 16'hB555, 16'hD619, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD619, 16'hD619, 16'hD619, 16'hD619, 16'hC596, 16'h5A89, 16'h9553, 16'h9D96, 16'h9D55, 16'h9D95, 16'h9D95, 16'h9D95, 16'hA5D6, 16'hA5D6, 16'h8512, 16'h9554, 16'h9D95, 16'h9D94, 16'h9D54, 16'h9D95, 16'h9D94, 16'h9D55, 16'h9D95, 16'h9D54, 16'h8CD2, 16'h9513, 16'h9D54, 16'h9D54, 16'h9D54, 16'h8CD1, 16'h634B, 16'h3000, 16'h6186, 16'hA451, 16'hD618, 16'hF71D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF1E, 16'hDD57, 16'hA24A, 16'h8800, 16'hA1C9, 16'hC2CD, 16'hCB8F, 16'hCC12, 16'hD493, 16'hBC52, 16'h5145, 16'h634B, 16'h6B4C, 16'h4186, 16'h7ACB, 16'hBD15, 16'hBD55, 16'h9C11, 16'h7B0C, 16'h4145, 16'h5B0B, 16'h8451, 16'h9D54, 16'hA5D5, 16'hA616, 16'h9553, 16'h5207, 16'hBDD6, 16'hFFDF, 16'hFFDF, 16'h8BCF, 16'h8CD2, 16'hA616, 16'hA5D6, 16'h9513, 16'h634B, 16'hD699, 16'hFF9E, 16'h9C51, 16'h7C0F, 16'h8C0F, 16'hF75D, 16'hFFDF, 16'hF75D, 16'h7B8D, 16'h9D94, 16'hAE57, 16'hAE57, 16'h9D54, 16'h52C9, 16'hBD95, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hD658, 16'hDE9A, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9C51, 16'h4042, 16'hC5D7, 16'hCE18, 16'h72CB, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'hC596, 16'hE6DB, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE18, 16'h8BCE, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h840F, 16'h9D54, 16'hAE17, 16'hAE17, 16'h8CD1, 16'h62CB, 16'h9513, 16'hAE17, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hA617, 16'hADD7, 16'h73CE, 16'h3986, 16'hB555, 16'hD619, 16'hD618,
        16'hD618, 16'hD618, 16'hD619, 16'hD619, 16'hD619, 16'hD618, 16'hD619, 16'h8B8F, 16'h740F, 16'hADD6, 16'h9D55, 16'h9D55, 16'h9D55, 16'h9D95, 16'h9D95, 16'h9D95, 16'h8D12, 16'h8D13, 16'hA5D6, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D54, 16'h9D95, 16'h9554, 16'h9513, 16'h9D54, 16'h9554, 16'h9554, 16'h9D95, 16'h9D94, 16'h9553, 16'h740F, 16'h4248, 16'h2000, 16'h6187, 16'h8B4E, 16'hBD15, 16'hEEDC, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hEE1A, 16'hB30E, 16'h9000, 16'hAA0A, 16'hC30E, 16'hCBD1, 16'hCC52, 16'hD493, 16'hCC92, 16'h9B0D, 16'h5145, 16'h2840, 16'h2000, 16'h000, 16'h40C3, 16'h730B, 16'h5A8A, 16'h4247, 16'h530B, 16'h4289, 16'h8491, 16'hA595, 16'hA595, 16'hA5D5, 16'hA5D6, 16'h8491, 16'h6289, 16'hD659, 16'hFFDF, 16'hFFDF,
        16'hC596, 16'h73CD, 16'hAE57, 16'hA595, 16'h740F, 16'h7B8D, 16'hDEDA, 16'hFFDF, 16'hDE9A, 16'h4985, 16'h9C92, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hB595, 16'h73CF, 16'hB658, 16'hA617, 16'h8491, 16'h5A89, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h72CB, 16'h730C, 16'hCE18, 16'h7B8E, 16'hBD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hE71C, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h7B0C, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB554, 16'h7C50, 16'hB617, 16'hB618, 16'h8CD2, 16'h9450, 16'h8C91, 16'hA5D6, 16'hAE17, 16'hADD6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hA617, 16'h8D13, 16'h5289, 16'h4186, 16'hAD14, 16'hD619, 16'hCE18, 16'hCE18, 16'hD619, 16'hD619, 16'hD619, 16'hD619, 16'hD619, 16'hB4D4, 16'h5249, 16'h9D54, 16'h9D95, 16'h9D95, 16'h9D55, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9553, 16'h7CD2, 16'h9DD6, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D55, 16'h9D95, 16'h9D54, 16'h9554, 16'h9554, 16'h9D54, 16'h9554, 16'h9554, 16'h9554, 16'h9D54, 16'h9D54, 16'h9D54, 16'h9513, 16'h7C4F, 16'h630B, 16'h3080, 16'h4800, 16'h7249, 16'hB4D3, 16'hD618,
        16'hEEDC, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF1E, 16'hEE19, 16'hCC11, 16'hA988, 16'hBA4B, 16'hCB8F, 16'hCC11, 16'hD493, 16'hD4D4, 16'hD4D4, 16'hD514, 16'hCCD4, 16'hC493, 16'hAB8F, 16'h5082, 16'h73CE, 16'h7C90, 16'h7C90, 16'h7C91, 16'h8D12, 16'h9D94, 16'h9554, 16'h638D, 16'h9D54, 16'hA595, 16'hA5D5, 16'h9D94, 16'h6BCE, 16'h834E, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h734C, 16'h9D94, 16'h84D1, 16'h630B, 16'hAD13, 16'hF79E, 16'hFFDF, 16'hF75D, 16'h9C51, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h734C, 16'hA596, 16'h9554, 16'h638C, 16'h8C0F, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h628A, 16'h7B8D, 16'hAD13, 16'h8B8E, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9C51, 16'hC5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDA, 16'h6B8C, 16'hAE16, 16'hB658, 16'h9513, 16'h9CD2, 16'hC5D6, 16'h7C50, 16'hB657, 16'hAE16,
        16'hADD6, 16'hADD6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'hAE17, 16'h9554, 16'h9491, 16'h6ACB, 16'h5289, 16'hA4D3, 16'hD618, 16'hCE18, 16'hCE18, 16'hD619, 16'hD619, 16'hD619, 16'hD619, 16'hD618, 16'h730B, 16'h740F, 16'hA5D6, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D94, 16'h7450, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D54, 16'h9D54, 16'h9554, 16'h9554, 16'h9D54, 16'h9554, 16'h9554, 16'h9554, 16'h9554, 16'h9554, 16'h9D95, 16'h8D12, 16'h8512, 16'hA5D5, 16'h9554, 16'h8CD1, 16'h73CE, 16'h4A47, 16'h4942, 16'h6186, 16'h8B8E, 16'hBD15, 16'hDE19, 16'hF71D, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF1D, 16'hEDD9, 16'hD412, 16'hC30D, 16'hC34F, 16'hCC11, 16'hD453, 16'hD494, 16'hD4D5, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hDD56, 16'hC452, 16'h50C2, 16'h8D12, 16'h9594, 16'h9594, 16'h9D94, 16'h9D94, 16'hA5D5,
        16'h7C50, 16'h73CE, 16'hA595, 16'h9D53, 16'h7C4F, 16'h730C, 16'hB555, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h6207, 16'h6B0B, 16'h7BCE, 16'hA4D2, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h730C, 16'h6B8D, 16'h7C0F, 16'h83CE, 16'hC617, 16'hFFDE, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h838E, 16'h730C, 16'h6ACB, 16'hCDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h8BCE, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h8C0F, 16'h8D13, 16'hB658, 16'hA595, 16'h7BCE, 16'hEF1C, 16'h9491, 16'h9553, 16'hB617, 16'hAE17, 16'hADD6, 16'hADD6, 16'hA617, 16'hAE17, 16'hA5D6, 16'hA5D6, 16'h9D95, 16'h8C91, 16'h8B8E, 16'hB555, 16'h9CD3, 16'h834D, 16'hCDD7, 16'hD619, 16'hCE18, 16'hCE18, 16'hD619, 16'hCE19, 16'hD619, 16'hBD55, 16'h4206, 16'h9D54, 16'hA595, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D95, 16'hA5D5, 16'h6C0F, 16'h8D13, 16'hA5D5, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D54, 16'h9D95, 16'h9554, 16'h84D2, 16'h9D94, 16'h9D54, 16'h9554,
        16'h9554, 16'h9554, 16'h9554, 16'h9D95, 16'h8CD2, 16'h744F, 16'h9594, 16'h9554, 16'h9594, 16'h9594, 16'h9D94, 16'h9D94, 16'h8CD1, 16'h73CE, 16'h4247, 16'h4100, 16'h5144, 16'h830D, 16'hAC92, 16'hCD96, 16'hEE9B, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5F, 16'hFF1D, 16'hEE5B, 16'hE556, 16'hD412, 16'hCBD1, 16'hD412, 16'hD494, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD556, 16'hBC51, 16'h4000, 16'h8CD1, 16'h9D95, 16'h9D95, 16'h9DD5, 16'h9594, 16'h744F, 16'h41C4, 16'h734D, 16'h7BCE, 16'h83CF, 16'hB555, 16'hEF1D, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hC5D7, 16'h8B8E, 16'hACD3, 16'hD659, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hC5D7, 16'h6ACA, 16'h838E, 16'hBD96, 16'hDEDB, 16'hFFDE, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hB514, 16'h4883, 16'h40C3, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9C50, 16'hCE18, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h6B8D, 16'hADD7, 16'hB617, 16'h638D, 16'hDEDA, 16'hEF1C, 16'h634C, 16'hA5D6, 16'hAE17, 16'hAE16, 16'hAE17, 16'hAE17, 16'hAE17, 16'hADD6, 16'hADD6, 16'hA5D6, 16'h84D1, 16'h734C, 16'hB555, 16'hEF5D, 16'h3944, 16'h5A48, 16'hA492, 16'hCDD7, 16'hD619, 16'hCE18, 16'hCE18, 16'hCE18, 16'hD619, 16'h93CF, 16'h5B0B, 16'hA595, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D95, 16'hA5D6, 16'h7C90, 16'h63CD, 16'hA5D6, 16'hA595, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D54, 16'h7C4F, 16'h9554, 16'h9D95, 16'h9554, 16'h9554, 16'h9554, 16'h9554, 16'h9D95, 16'h8CD2, 16'h6BCD, 16'h9D95, 16'h9594, 16'h9553, 16'h9553, 16'h8D53, 16'h8D53, 16'h9593, 16'h9593, 16'h9594, 16'h8D12, 16'h740E, 16'h634B, 16'h4A47, 16'h2880, 16'h4000, 16'h728A, 16'h9BCF, 16'hBC93, 16'hCD56, 16'hD597, 16'hDDD8, 16'hE5D8, 16'hDD56, 16'hD493, 16'hCBD1, 16'hCB90, 16'hCBD1, 16'hD453, 16'hD4D4, 16'hD4D5, 16'hD4D5, 16'hD4D5, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515,
        16'hD515, 16'hD515, 16'hD515, 16'hDD56, 16'hBC11, 16'h4103, 16'h8CD2, 16'h8CD2, 16'h7C50, 16'h6BCE, 16'h630B, 16'hA4D3, 16'hC5D7, 16'hCE17, 16'hE6DB, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hEF1C, 16'hFFDE, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hD699, 16'hCE18, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DA, 16'h8BCF, 16'h6208, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hA410, 16'hF75C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDE, 16'h8C50, 16'h9513, 16'hBE58, 16'h8491, 16'hAD54, 16'hFFDF, 16'hC617, 16'h638C, 16'hAE17, 16'hAE17, 16'hAE17, 16'hAE17, 16'hAE17, 16'hADD6, 16'hADD6, 16'hAE17, 16'h8D13, 16'h7C0E, 16'h8C0E, 16'hFF9E, 16'hA4D3, 16'h634C, 16'h738D, 16'h730B, 16'hA492, 16'hC596, 16'hD619, 16'hD619, 16'hD619, 16'hCDD7, 16'h6289, 16'h7C50, 16'hA5D6, 16'h9D95, 16'h9DD5, 16'h9D95, 16'hA5D6, 16'h8D13, 16'h4AC8, 16'h7C4F,
        16'hADD6, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D95, 16'hA595, 16'h8490, 16'h7C4F, 16'h9D94, 16'h9554, 16'h9554, 16'h9554, 16'h9554, 16'h9D95, 16'h8CD2, 16'h4246, 16'h8D12, 16'h9D95, 16'h9554, 16'h8D12, 16'h8D53, 16'h8D53, 16'h8D53, 16'h8D53, 16'h8D53, 16'h8511, 16'h7490, 16'h8D53, 16'h9553, 16'h8D12, 16'h8C91, 16'h5A8A, 16'h1800, 16'h6000, 16'h6000, 16'h7800, 16'h9803, 16'hB1C9, 16'hBA8C, 16'hC34F, 16'hCBD1, 16'hD454, 16'hD4D5, 16'hD4D5, 16'hD4D5, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD556, 16'hBC52, 16'h2800, 16'h62CB, 16'h8C10, 16'hA4D3, 16'hCE18, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE18, 16'h9C50, 16'hD659, 16'hFF9E,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'hBD54, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h6BCD, 16'hB657, 16'hA595, 16'h840F, 16'hF79E, 16'hFFDF, 16'hAD14, 16'h6BCD, 16'hAE17, 16'hAE17, 16'hAE17, 16'hAE17, 16'hADD7, 16'hADD7, 16'hAE17, 16'h9D95, 16'h7C50, 16'h62CA, 16'hEF1C, 16'hD659, 16'h634C, 16'hB658, 16'h9D54, 16'h5289, 16'h5208, 16'h8BCF, 16'hC596, 16'hD618, 16'hD619, 16'hBD55, 16'h4A07, 16'h8D12, 16'hA5D6, 16'h9DD5, 16'hA5D6, 16'hA5D6, 16'h9594, 16'h9490, 16'h940F, 16'h7C4F, 16'hA5D6, 16'h9D96, 16'hA595, 16'hA595, 16'hA595, 16'h9D95, 16'hA596, 16'h9513, 16'h4246, 16'h8CD1, 16'h9D95, 16'h9554, 16'h9D95, 16'h9D54, 16'h9D95, 16'h84D2, 16'h9491, 16'h738D, 16'h9554, 16'h9D95, 16'h7C91, 16'h5B8C, 16'h8D53, 16'h8D53, 16'h8D53, 16'h8D53, 16'h8512, 16'h5BCD, 16'h8512, 16'h8512, 16'h8512, 16'h8552, 16'h8CD1, 16'h59C7, 16'h9209, 16'hAA4A, 16'hAA8B, 16'hBB0E, 16'hCB90, 16'hCC12, 16'hD493, 16'hD4D5, 16'hD4D5,
        16'hD4D5, 16'hD4D5, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD516, 16'hD515, 16'hDD56, 16'hBC52, 16'h3800, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hEF5C, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9C91, 16'h8CD1, 16'hBE58, 16'h738D, 16'hD659, 16'hFFDF, 16'hFF9E, 16'h9CD2, 16'h6BCD, 16'hA617, 16'hB658, 16'hAE17, 16'hAE17, 16'hAE17, 16'hAE17, 16'hAE16, 16'h7C51, 16'h5ACA, 16'hC5D7, 16'hFF9E, 16'h5A89, 16'h9D54, 16'hBE99, 16'h8491, 16'h8C50, 16'hB554, 16'h51C5,
        16'h7B4D, 16'hACD3, 16'hD5D7, 16'hB4D3, 16'h5ACA, 16'h9514, 16'hA617, 16'hA5D6, 16'hA5D6, 16'h9DD6, 16'h844F, 16'hDE99, 16'hA4D3, 16'h740E, 16'hA5D6, 16'hA5D6, 16'hA595, 16'h9D95, 16'h9D95, 16'h9D95, 16'h9D95, 16'h7C0E, 16'h73CD, 16'h9512, 16'h9D95, 16'h9554, 16'h9D95, 16'h9DD5, 16'h744F, 16'hDEDA, 16'hC617, 16'h634B, 16'hA616, 16'h8D12, 16'h4287, 16'h5B8B, 16'h8D12, 16'h9594, 16'h8D93, 16'h8D94, 16'h6C4F, 16'h7490, 16'h8D53, 16'h8512, 16'h8512, 16'h8D12, 16'h5249, 16'h7146, 16'hCBD1, 16'hC411, 16'hCC53, 16'hD494, 16'hD4D5, 16'hD4D5, 16'hD4D5, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD516, 16'hD516, 16'hD515, 16'hDD56, 16'hBC52, 16'h4000, 16'hD617, 16'hDE9A, 16'hDE59, 16'hDE59, 16'hDE59, 16'hE6DB, 16'hEF1B, 16'hF75D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5C, 16'h734C, 16'h9D13, 16'h9513, 16'h9451, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB555, 16'h6B8D, 16'h9D95, 16'hB658, 16'hAE17, 16'hAE17, 16'hAE17, 16'hAE57, 16'h9553, 16'h5B0B, 16'h9C51, 16'hFFDF, 16'hBD96, 16'h5ACA, 16'hB658, 16'hA595, 16'h8450, 16'hFFDF, 16'hCE18, 16'h800, 16'h5ACA, 16'h6ACA, 16'h8BCE, 16'h5A08, 16'h3985, 16'h7C50, 16'h9554, 16'h9DD5, 16'hAE57, 16'h7C90, 16'hB554, 16'hFFDF, 16'hACD3, 16'h638C, 16'h9D54, 16'hAE17, 16'hA5D6, 16'hA5D6, 16'h9D95, 16'hA596, 16'h8C91, 16'hAD13, 16'h7BCE, 16'h84D1, 16'h9D95, 16'h9594, 16'hA5D6, 16'h744F, 16'hD69A, 16'hFFDF, 16'hA4D2, 16'h6BCD, 16'h9553, 16'hA554, 16'hCE58, 16'h5B4A, 16'h6C8F, 16'h8552, 16'h9594, 16'h8D53, 16'h32C8, 16'h8D53, 16'h9594,
        16'h8D53, 16'h9D94, 16'h9451, 16'h4800, 16'hCC93, 16'hD4D5, 16'hD4D5, 16'hD4D5, 16'hD4D5, 16'hD4D5, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hDD56, 16'hBC52, 16'h4800, 16'h5144, 16'h4944, 16'h4945, 16'h5144, 16'h4881, 16'h5945, 16'h61C7, 16'h6208, 16'h830D, 16'hBD14, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h628A, 16'h8491, 16'h7BCE, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h738D, 16'h84D2, 16'hAE57, 16'hB658, 16'hAE17,
        16'hAE17, 16'hAE17, 16'h7C50, 16'h5A88, 16'hE6DB, 16'hFFDF, 16'h7B4D, 16'h8CD2, 16'hBE59, 16'h73CE, 16'hCE17, 16'hFFDF, 16'hC5D7, 16'h6B8E, 16'h9554, 16'h8CD2, 16'h7C50, 16'h7C50, 16'h52C9, 16'h7C90, 16'hA616, 16'hAE57, 16'hA5D6, 16'h6B8C, 16'hEF5C, 16'hFFDF, 16'hCE18, 16'h7BCD, 16'h744F, 16'h9D94, 16'hA5D6, 16'hA5D6, 16'hA5D6, 16'h9D55, 16'h8C10, 16'hD659, 16'h7BCE, 16'h7C90, 16'hA5D6, 16'hAE17, 16'h7C4F, 16'hD699, 16'hFFDF, 16'hFFDF, 16'hC5D7, 16'h630A, 16'h8C10, 16'hFFDF, 16'hF79E, 16'hC5D7, 16'h8C51, 16'h73CE, 16'h7C0F, 16'hA513, 16'h73CD, 16'h7C50, 16'h7C4F, 16'h844F, 16'h730B, 16'h3800, 16'hC452, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD516, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD556, 16'hC493, 16'h4000, 16'h83CE, 16'h9D13, 16'h9D13, 16'h9D13, 16'hA513, 16'hA554, 16'hA554, 16'hA513, 16'h9CD2, 16'h4986, 16'h834D, 16'hFF9E, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h7B4D, 16'h5A89, 16'h62CA, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h9C91, 16'h6B8D, 16'h9553, 16'hAE17, 16'hAE58, 16'hB658, 16'hA5D6, 16'h5B4C, 16'h9450, 16'hFFDF, 16'hDE9A, 16'h5248, 16'hB617, 16'hADD6, 16'h7B8D, 16'hF79E, 16'hFFDF, 16'hCE18, 16'h7BCF, 16'hA595, 16'hB699, 16'hB698, 16'h9D95, 16'h5B4C, 16'h9513, 16'hB658, 16'hB698, 16'h8491, 16'hA4D3, 16'hFFDF, 16'hFFDF, 16'hF79D, 16'hBD95, 16'h738D, 16'h6BCE, 16'h8D13, 16'hA5D6, 16'hB617, 16'h9513, 16'h9C92, 16'hEF1C, 16'hA493, 16'h6BCD, 16'hAE16, 16'h7C90, 16'hD699, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hEF1C, 16'h8BCF, 16'hB555, 16'hCE18, 16'hBD95, 16'h8B8E, 16'h4000, 16'h4903, 16'h9410, 16'h5A08, 16'h5A48, 16'h8C10, 16'h9CD3, 16'hACD3, 16'h4903, 16'hA38F, 16'hD516, 16'hD4D5, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD516, 16'hD515, 16'hD516, 16'hD516, 16'hD555, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD516, 16'hCCD4, 16'h58C4, 16'h6B4C, 16'h9D13, 16'h9512, 16'h9D53, 16'hA554, 16'h9491, 16'h7BCD, 16'hB5D5, 16'hCE99, 16'hC617, 16'h000, 16'hC5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hF79E, 16'hAD14, 16'h3040, 16'h5207, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h8C10, 16'h634C, 16'h6C0E, 16'h84D2, 16'h9D95, 16'h9D94, 16'h4248, 16'hC5D7, 16'hFFDF, 16'hBD95, 16'h6B8D, 16'hBE99, 16'h8490, 16'hAD14, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h8C0F, 16'h7C90, 16'hA616, 16'hB699, 16'hA616, 16'h638D, 16'h7C90, 16'hAE58, 16'hBE98, 16'h73CE, 16'hCE58, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hCE18, 16'h9450, 16'h738D, 16'h740F, 16'h9513, 16'h5B0A, 16'h8C10, 16'hE71C, 16'hBD96, 16'h840F, 16'h5309, 16'hD699, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h8BCF, 16'h6ACA, 16'h6249, 16'h730B, 16'h83CE, 16'h9450, 16'hA513, 16'hAD55, 16'hAD95, 16'hBDD6, 16'hC618, 16'hC658, 16'hC659, 16'hC617, 16'h4944, 16'h9B4E, 16'hD516, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD516, 16'hD516, 16'hD516, 16'hD515, 16'hD516, 16'hD556, 16'hD516, 16'hD516, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD516, 16'hD4D4, 16'h79C7, 16'h5207, 16'h9CD2,
        16'hA554, 16'h9CD2, 16'h6B0B, 16'h4183, 16'h9CD2, 16'hC658, 16'hC618, 16'hCE58, 16'h7B8D, 16'h838E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71D, 16'hD6DB, 16'hD6DC, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h9450, 16'h72CA, 16'hD618, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'hB595, 16'h8C50, 16'h7B8D, 16'h7BCE, 16'h6B0C, 16'h59C6, 16'hDE9A, 16'hFFDF, 16'h9C50, 16'h6BCE, 16'hBE18, 16'h7BCE, 16'hCE58, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hAD14, 16'h6B4C, 16'h8CD2, 16'hAE17, 16'hBE58, 16'h8491, 16'h6BCD, 16'h9D54, 16'hADD6, 16'h734C, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hEF1C, 16'hCE18, 16'hBD95, 16'hAD54, 16'h9451, 16'h9C91, 16'hE71B, 16'hFF9E, 16'hACD3, 16'hB555, 16'hFFDF, 16'hFFDF, 16'hA492, 16'h41C6, 16'hC617, 16'hCE59, 16'hCE99, 16'hCE9A, 16'hCE99, 16'hC659, 16'hC658, 16'hC658, 16'hC658, 16'hBE18, 16'hBE17, 16'hBE17, 16'hC618, 16'h730C, 16'h8ACC, 16'hD515, 16'hCD15, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD516, 16'hD516, 16'hD555, 16'hD515, 16'hD515, 16'hD516, 16'hD516, 16'hD515, 16'hD516, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hB3D0, 16'h4000, 16'h730B, 16'h838E, 16'h40C2, 16'h6ACB, 16'hB595, 16'hC658, 16'hC618, 16'hC618, 16'hCE59, 16'h9C92, 16'h59C7, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE75D, 16'hC65A, 16'hCE9B, 16'hC65A, 16'hD6DC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'hCE18, 16'hDEDA, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hEF1C, 16'hEF5C, 16'hDEDA, 16'hA4D2, 16'hE71C, 16'hFF9E, 16'h9C91, 16'h6B0C, 16'h9492, 16'h62CA, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'hACD3, 16'h8C0F, 16'h9D12, 16'hBDD6, 16'hC618, 16'hAD13, 16'h9491, 16'h738D, 16'h4143, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hFFDF, 16'hF75D, 16'h3800, 16'hB5D6, 16'hCE99, 16'hBE17, 16'hAD95, 16'hAD95, 16'hB5D6, 16'hC658, 16'hC658, 16'hC618, 16'hBE17, 16'hBE17, 16'hB5D6, 16'hAD54, 16'hAD54, 16'h5A49, 16'h8ACB, 16'hD515, 16'hCD15, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515,
        16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hCD15, 16'hD515, 16'hD556, 16'hD514, 16'h7A08, 16'h000, 16'h5A08, 16'hA4D3, 16'hCE18, 16'hCE58, 16'hC658, 16'hC658, 16'hC658, 16'hCE59, 16'hB595, 16'h3800, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD6DB, 16'hCE9B, 16'hDF1D, 16'hD69B, 16'hCE9B, 16'hF79F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hD658, 16'h9C91, 16'h6B0B, 16'h000, 16'h8BCF, 16'hD699, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hF75D,
        16'hE6DB, 16'hDEDB, 16'hFF9E, 16'hFFDF, 16'hF75D, 16'hDEDB, 16'hC5D7, 16'h9C10, 16'hBD55, 16'hEF1D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD56, 16'h6B0B, 16'hCE99, 16'hCE99, 16'h9D13, 16'h7BCD, 16'h8C8F, 16'h8C4F, 16'h9CD2, 16'hA553, 16'hAD54, 16'h9CD2, 16'h9491, 16'h8C90, 16'h844F, 16'h8C4F, 16'h41C6, 16'h828B, 16'hDD15, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD516, 16'hD516, 16'hD515, 16'hD515, 16'hD515, 16'hD516, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD556, 16'hDD56, 16'hD515, 16'hB410, 16'h69C7, 16'h4944, 16'h9410, 16'hCE18, 16'hCE59, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hCE59, 16'hC618, 16'h3882, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hDEDB, 16'hCE18, 16'hAD14, 16'hAD14, 16'hA4D3, 16'hA492, 16'hC597, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE75D, 16'hC69A, 16'hDF1C, 16'hF7DF, 16'hD69B, 16'hCE9B, 16'hF7DF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5C, 16'hD658, 16'hAD14, 16'hAD13, 16'hC5D7, 16'hE6DA, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hF79D, 16'hFFDF, 16'hFF9F, 16'hE6DB, 16'hB596, 16'h9C51, 16'h838E, 16'h7B0D, 16'hDE9B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h7B4E, 16'h9CD2, 16'hCE99, 16'hC659, 16'hA513, 16'h2000, 16'h840F, 16'h9490, 16'h844F, 16'h840F, 16'h844F, 16'h844F, 16'h8C4F, 16'h8C90, 16'h8C90, 16'h9490, 16'h5248, 16'h828B, 16'hD515, 16'hCD15, 16'hD515,
        16'hD515, 16'hD516, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hCD15, 16'hD515, 16'hD556, 16'hDD56, 16'hCCD4, 16'hA38F, 16'h6986, 16'h5A08, 16'h9451, 16'hC5D7, 16'hCE58, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hCE59, 16'h5249, 16'hB554, 16'hFFDF, 16'hE6DB, 16'hC597, 16'h9410, 16'h8B8F, 16'h6A4A, 16'h72CB, 16'h830C, 16'h8B8E, 16'h8B4D, 16'h834D, 16'h8B8F, 16'h5145, 16'h5146, 16'hC596, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD6DC,
        16'hC69A, 16'hF79E, 16'hEF5E, 16'hC65A, 16'hD6DC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE75D, 16'hD69B, 16'hD6DC, 16'hEF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hCDD7, 16'h728A, 16'h2800, 16'h6289, 16'h83CE, 16'hA492, 16'h8BCF, 16'h5A07, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h6249, 16'hB5D6, 16'hC659, 16'hC618, 16'hCE58, 16'h9C92, 16'h3081, 16'h840E, 16'h9490, 16'h8C90, 16'h8C90, 16'h8C50, 16'h8C90, 16'h8C90, 16'h8C90, 16'h8C4F, 16'h4144, 16'h92CC, 16'hD515, 16'hCD15, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD556, 16'hD515, 16'hD515, 16'hCD15, 16'hD515, 16'hD515, 16'hD515, 16'hCD15, 16'hD556, 16'hD556, 16'hD556, 16'hC493, 16'h930C, 16'h6186, 16'h72CB, 16'hB4D4, 16'hCE18, 16'hD659, 16'hCE59, 16'hC618, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hCE59, 16'h7BCF, 16'h3882, 16'h938E, 16'h5143, 16'h5185, 16'h9C51, 16'hB4D3, 16'hC596, 16'hC596, 16'hBD96, 16'hBD55,
        16'h93CF, 16'hA492, 16'hD618, 16'hC618, 16'hA4D3, 16'h3800, 16'h7ACC, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5E, 16'hC69B, 16'hD6DC, 16'hFFDF, 16'hE71D, 16'hC69B, 16'hDF1D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79F,
        16'hCE9B, 16'hCE9B, 16'hC69B, 16'hCE9B, 16'hEF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'hA492, 16'h59C8, 16'h5145, 16'h9451, 16'hB596, 16'hC658, 16'hCE58, 16'hCE99, 16'hCE58, 16'h940F, 16'h3000, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h4144, 16'hC618, 16'hC658, 16'hC618, 16'hC618, 16'hCE59, 16'hA4D3, 16'h2800, 16'h7B8D,
        16'h9490, 16'h8C90, 16'h8C90, 16'h8C90, 16'h8C90, 16'h8C91, 16'h840F, 16'h2800, 16'h930D, 16'hD515, 16'hD515, 16'hD515, 16'hCD15, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD516, 16'hD515, 16'hD515, 16'hCD15, 16'hCD15, 16'hD516, 16'hD556, 16'hD514, 16'hABCF, 16'h7208, 16'h5946, 16'h838E, 16'hBD56, 16'hD619, 16'hD659, 16'hCE58, 16'hCE58, 16'hCE58, 16'hC658, 16'hC618, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC618, 16'hCE59, 16'hA513, 16'h38C2, 16'hAC92, 16'h93CF, 16'hB514, 16'hC5D7, 16'hB554, 16'hAD14, 16'hA4D2, 16'hA4D3, 16'h9410, 16'h7B0C, 16'hBD95, 16'hC617, 16'hC618, 16'hCE58, 16'hBD96, 16'h83CE, 16'h3800, 16'hB514, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDC, 16'hC65A, 16'hE71D, 16'hFFDF, 16'hD6DC, 16'hCE9B, 16'hEF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hCE9B, 16'hD6DC, 16'hDF1D, 16'hCE9B, 16'hCE9B, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hACD3, 16'h2800, 16'h6289, 16'hA4D3, 16'hC617, 16'hCE58, 16'hC618, 16'hBDD7, 16'hBD96, 16'hBD96, 16'h8C0F, 16'h8B8D, 16'h9C51, 16'h4145, 16'hC5D7, 16'hFF9E, 16'hB4D4, 16'h630B, 16'hCE59, 16'hC618, 16'hC658, 16'hC658, 16'hC658, 16'hCE59, 16'hA4D2, 16'h800, 16'h7B4D, 16'h94D1, 16'h8C90, 16'h8C91, 16'h8C90, 16'h94D1, 16'h83CE, 16'h000, 16'h9B4E, 16'hD516, 16'hCD15, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hCD15, 16'hD556, 16'hDD56, 16'hD515, 16'hC493, 16'h930D, 16'h5104, 16'h6A89, 16'h9C50, 16'hC597, 16'hD659, 16'hCE59, 16'hC618, 16'hCE59, 16'hCE58, 16'hCE58, 16'hC658, 16'hCE58, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658,
        16'hCE59, 16'hB555, 16'h51C7, 16'hA451, 16'h838D, 16'hAD14, 16'hA513, 16'hAD13, 16'hA4D3, 16'hA4D3, 16'hA492, 16'h72CB, 16'h9C51, 16'hAD14, 16'hBE17, 16'hC618, 16'hC618, 16'hC658, 16'hCE58, 16'hAD14, 16'h4843, 16'h8B8E, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69B, 16'hCE9B, 16'hF79E, 16'hF79F, 16'hCE9B, 16'hD69B, 16'hF79F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79F, 16'hCE9B, 16'hD6DC, 16'hF7DF, 16'hD6DC, 16'hC65A, 16'hDEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE18, 16'h5145, 16'h5A49, 16'hAD54, 16'hCE58, 16'hC658, 16'hBE17, 16'hBE17, 16'hBDD7, 16'hBDD6, 16'h9450, 16'h9450, 16'h9C51, 16'h9451, 16'hBDD6, 16'hA451,
        16'h2800, 16'h59C8, 16'h3842, 16'h94D2, 16'hCE99, 16'hC618, 16'hC658, 16'hC658, 16'hC618, 16'hC618, 16'hCE59, 16'hA4D3, 16'h3000, 16'h734C, 16'h94D1, 16'h94D1, 16'h94D1, 16'h9491, 16'h49C7, 16'h5000, 16'hAB90, 16'hD516, 16'hCD15, 16'hD515, 16'hD515, 16'hCD15, 16'hD515, 16'hD556, 16'hD556, 16'hDD56, 16'hD515, 16'hC493, 16'h9B8E, 16'h7208, 16'h5945, 16'h838E, 16'hB555, 16'hD659, 16'hD659, 16'hD659, 16'hCE58, 16'hC618, 16'hCE59, 16'hCE59, 16'hCE58, 16'hCE59, 16'hC658, 16'hCE58, 16'hCE59, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC617, 16'h5248, 16'h59C6, 16'hA492, 16'hAD14, 16'hAD14, 16'hAD14, 16'hAD13, 16'hB555, 16'h9410, 16'h5A08, 16'h9C51, 16'hB554, 16'hC617, 16'hC618, 16'hC618, 16'hC618, 16'hC618, 16'hC618, 16'hC5D6, 16'h6249, 16'h830C, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF9E, 16'hCE9B, 16'hD6DB, 16'hFFDF, 16'hE71D, 16'hC69B, 16'hDF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD6DC, 16'hC65A, 16'hF79F, 16'hEF9E, 16'hCE9B, 16'hCE9B, 16'hEF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h9C51, 16'h2800, 16'h9C91, 16'hCE58, 16'hCE99, 16'hCE99, 16'hCE99, 16'hC658, 16'hC618, 16'hC617, 16'hBD96, 16'h838D, 16'hA4D3, 16'hBDD6, 16'hB5D6, 16'hBDD6, 16'hA492, 16'hA451, 16'h8C0F, 16'h000, 16'hB595, 16'hCE99, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC618, 16'hC658, 16'hCE59, 16'hB555, 16'h4104, 16'h6B4B, 16'h9D12, 16'h9CD2, 16'h6ACA, 16'h6946, 16'hB30E, 16'hC493, 16'hD515, 16'hCD15, 16'hCD15, 16'hD515, 16'hD556, 16'hDD56, 16'hD515, 16'hBC52, 16'h9B4E, 16'h7209, 16'h61C7, 16'h7B4D, 16'hA4D3, 16'hC5D7, 16'hD659, 16'hD699, 16'hCE59, 16'hCE58, 16'hCE58, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE58,
        16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hC658, 16'hC658, 16'hCE58, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hCE59, 16'h734D, 16'h4985, 16'hB514, 16'hAD14, 16'hAD13, 16'hAD54, 16'hB554, 16'h9450, 16'h3080, 16'h730C, 16'hBD55, 16'hC618, 16'hC618, 16'hC618, 16'hC618, 16'hC618, 16'hC618, 16'hC618, 16'hC618, 16'hC618, 16'h6A8A, 16'h72CB, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5E, 16'hC65A, 16'hDF1D, 16'hFFDF, 16'hD69B, 16'hCE9B, 16'hEF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71D, 16'hC65A, 16'hE71D, 16'hFFDF, 16'hE71C, 16'hC69B, 16'hD6DC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h72CB, 16'h5186, 16'hBDD6, 16'hCE99, 16'hC617, 16'hBD96,
        16'hB595, 16'hAD54, 16'hB555, 16'hBDD6, 16'hBDD7, 16'hAD14, 16'h83CF, 16'hB595, 16'hB596, 16'hB596, 16'hB596, 16'hAD13, 16'h944F, 16'h9C91, 16'h2944, 16'hBE17, 16'hCE59, 16'hC658, 16'hC658, 16'hC618, 16'hC618, 16'hC618, 16'hC618, 16'hC658, 16'hCE59, 16'hBD96, 16'h5A49, 16'h62CA, 16'h730C, 16'h48C3, 16'hB411, 16'hCD15, 16'hCD15, 16'hCD15, 16'hD556, 16'hD556, 16'hD515, 16'hBC52, 16'h930C, 16'h7207, 16'h6249, 16'h83CF, 16'hAD14, 16'hC617, 16'hD659, 16'hD69A, 16'hCE59, 16'hCE58, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hC658, 16'hC658, 16'hC658, 16'hCE58, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hCE59, 16'h9491, 16'h2800, 16'hB514, 16'hBD96, 16'hBD96, 16'hACD3, 16'h6A8A, 16'h48C2, 16'h9410, 16'hCE18, 16'hCE59, 16'hCE58, 16'hCE58, 16'hC618, 16'hC658, 16'hC618, 16'hC617, 16'hC618, 16'hC617, 16'hC617, 16'hC5D7, 16'h624A, 16'h8B8E, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5E, 16'hCE9B, 16'hDEDC, 16'hDF1C, 16'hCE9B, 16'hD6DC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79F, 16'hCE9B, 16'hCE9B, 16'hF79F, 16'hF79F, 16'hCE9B, 16'hCE9B, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h6209, 16'h730C, 16'hCE58, 16'hC658, 16'hA514, 16'h83CE, 16'h9C51, 16'hA492, 16'h9C51, 16'h9C51, 16'hAD54, 16'hA513, 16'h734C, 16'h9CD2, 16'hB596, 16'hB596, 16'hB596, 16'hB595, 16'hB595, 16'hA4D2, 16'h730B, 16'h630B, 16'hCE58, 16'hC658, 16'hC658, 16'hC618, 16'hC618, 16'hC618, 16'hC618, 16'hC618, 16'hC658, 16'hC618, 16'hCE59, 16'hC5D7, 16'h734D, 16'h2000, 16'hB452, 16'hD556, 16'hCD15, 16'hCD15, 16'hD556, 16'hCCD4, 16'h930D, 16'h69C6, 16'h7B0B, 16'h9C91, 16'hBD96, 16'hD659, 16'hD699, 16'hD699, 16'hCE59,
        16'hC658, 16'hCE58, 16'hCE58, 16'hCE59, 16'hCE58, 16'hCE58, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hCE59, 16'hA513, 16'h000, 16'h6B0B, 16'hACD3, 16'h9C50, 16'h2800, 16'h6A8A, 16'hA492, 16'hACD4, 16'hBD96, 16'hCE18, 16'hCE58, 16'hCE58, 16'hC618, 16'hCE58, 16'hC618, 16'hC618, 16'hC618, 16'hC618, 16'hC5D7, 16'hC618, 16'hBD96, 16'h2000, 16'hBD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79F, 16'hCE9B, 16'hCE9B, 16'hCE9B, 16'hCE9B, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDC, 16'hC65A, 16'hE71D, 16'hFFDF, 16'hDEDC, 16'hC65A, 16'hE75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC597, 16'h6248, 16'hCE58, 16'hB595, 16'h8C10, 16'h9451, 16'hB556, 16'hCE18, 16'hCE18, 16'hCE18, 16'hCE18, 16'hC618, 16'hAD14, 16'h5A08, 16'hAD14, 16'hAD95, 16'hB595, 16'hB595, 16'hBD96, 16'hBD95, 16'hB554, 16'h3103, 16'h8410, 16'hCE59, 16'hC618, 16'hC618, 16'hC618, 16'hC658, 16'hC618, 16'hC618, 16'hC618, 16'hC658, 16'hC658, 16'hC658, 16'hCE58, 16'hCE18, 16'h9410, 16'h4883, 16'hB410, 16'hD515, 16'hCD15, 16'hBC52, 16'h69C7, 16'h9C92, 16'hCE59, 16'hDE9A, 16'hD69A, 16'hD659, 16'hC659, 16'hC658, 16'hCE58, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE58, 16'hCE58, 16'hCE59, 16'hCE59, 16'hCE59, 16'hC658, 16'hCE58, 16'hCE59, 16'hC658, 16'hCE58, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hCE59, 16'hC618, 16'h9CD2, 16'h9450, 16'h62CA, 16'h000, 16'h3000, 16'h9410, 16'hCDD8, 16'hC5D7, 16'hACD3, 16'h9C92, 16'hACD3, 16'hC5D7, 16'hCE59, 16'hCE58, 16'hC618, 16'hC618, 16'hC618, 16'hC618,
        16'hC617, 16'hC618, 16'hC618, 16'hC618, 16'h9C51, 16'h5145, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5E, 16'hD6DC, 16'hDEDC, 16'hEF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5E, 16'hC65B, 16'hCE9B, 16'hFFDF, 16'hEF5E, 16'hC65A, 16'hDF1C,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hEF1C, 16'hDE9A, 16'hC596, 16'h5A08, 16'h9C51, 16'hB555, 16'h7B0C, 16'hACD3, 16'hCE18, 16'hC618, 16'hCE18, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE59, 16'hBD96, 16'h5A08, 16'hA4D3, 16'hB595, 16'hB595, 16'hBD95, 16'h9410, 16'h5249, 16'h49C6, 16'h000, 16'h9D13, 16'hCE59, 16'hC658, 16'hC658, 16'hC618, 16'hC658, 16'hC658, 16'hC658, 16'hC618, 16'hC618, 16'hC658, 16'hCE58, 16'hC658, 16'hCE58, 16'hD699, 16'hAD14, 16'h4000, 16'hABCF,
        16'hC4D3, 16'h5986, 16'h9C51, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hEF5D, 16'hE71C, 16'hD69A, 16'hD659, 16'hCE59, 16'hCE59, 16'hC618, 16'hCE58, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE58, 16'hCE59, 16'hCE59, 16'hCE58, 16'hCE59, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE59, 16'hCE58, 16'hCE59, 16'hCE59, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE59, 16'hC658, 16'hCE59, 16'hAD54, 16'h9C91, 16'hA4D2, 16'h6248, 16'h4986, 16'hB514, 16'hD659, 16'hCE19, 16'hD619, 16'hCE18, 16'hBD56, 16'hA492, 16'hA493, 16'hC5D6, 16'hCE59, 16'hCE18, 16'hC618, 16'hC618, 16'hC618, 16'hC618, 16'hC618, 16'hC618, 16'hC618, 16'hBDD6, 16'h3000, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD6DC, 16'hC65A, 16'hE75D, 16'hF79E, 16'hC69B, 16'hD6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hDE9A, 16'hC596, 16'h9C50, 16'h728A, 16'h4080, 16'h2000, 16'h38C3, 16'h4104, 16'h8BCF, 16'h8BCF, 16'hB555, 16'hC618, 16'hC618, 16'hCE18, 16'hD659, 16'hCE59, 16'hCE58, 16'hCE59, 16'hCE59, 16'hCE59, 16'h7B0D, 16'h8BCF, 16'hB595, 16'hBD96, 16'h8BCE, 16'h1800, 16'h6B4C, 16'h8C50, 16'h3104, 16'hB596, 16'hCE59, 16'hC658, 16'hC658, 16'hCE58, 16'hC618, 16'hC618, 16'hC618, 16'hC618, 16'hC658, 16'hC658, 16'hC658, 16'hCE59, 16'hC618, 16'h8C0F, 16'h8BCF, 16'h8B8E, 16'h6208, 16'h7208, 16'h7B4D, 16'h83CE, 16'h4186, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hF79E, 16'hEF5D, 16'hE71C, 16'hDEDB, 16'hDE9A, 16'hD69A, 16'hCE99, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE59, 16'hD69A, 16'hD69A, 16'hCE59, 16'hCE58, 16'hCE59, 16'hCE59, 16'hCE58, 16'hCE59, 16'hCE59, 16'hC658, 16'hCE59, 16'hCE59, 16'hBDD6, 16'hA512, 16'h83CE, 16'h3800, 16'h7B4C, 16'hC5D7, 16'hD659, 16'hCE18,
        16'hCE19, 16'hCE18, 16'hCE19, 16'hCE19, 16'hBD96, 16'hA492, 16'hA492, 16'hC5D7, 16'hCE18, 16'hC618, 16'hC618, 16'hC618, 16'hC618, 16'hC617, 16'hC618, 16'hC618, 16'hCE58, 16'h730C, 16'h940F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5E, 16'hC65A, 16'hD6DB, 16'hD6DC, 16'hC65A, 16'hD6DC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'hAD13, 16'h7B4D, 16'h5145, 16'h40C2, 16'h5A49, 16'h838E, 16'h9C92, 16'hAD14, 16'hC5D7, 16'hBD55, 16'h4083, 16'h834E, 16'hBD96, 16'hCE18, 16'hC618, 16'hCE18, 16'hCE19, 16'hCE59, 16'hD659, 16'hD659, 16'hCE18, 16'hC596, 16'hC5D7, 16'h9410, 16'h6A8A, 16'hBD96, 16'h9C10, 16'h3882, 16'h94D2, 16'hBDD6, 16'h734C, 16'h62CA, 16'hC618, 16'hC658, 16'hC618, 16'hC618, 16'hC618, 16'hCE58,
        16'hCE58, 16'hC658, 16'hCE58, 16'hCE59, 16'hC658, 16'hC618, 16'hD659, 16'h8C0F, 16'h6ACB, 16'hA492, 16'h734D, 16'h30C2, 16'h000, 16'hA4D2, 16'hA514, 16'h5A89, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hF79E, 16'hF79E, 16'hF79D, 16'hF79D, 16'hF79E, 16'hF79E, 16'hF79E, 16'hFF9E, 16'hDEDA, 16'hCE58, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE58, 16'hCE59, 16'hCE59, 16'hC658, 16'hC617, 16'hAD13, 16'h6ACB, 16'h4145, 16'hACD3, 16'hD619, 16'hD659, 16'hCE19, 16'hCE19, 16'hCE19, 16'hCE18, 16'hCE18, 16'hCE18, 16'hCE59, 16'hBD96, 16'hA492, 16'hA4D3, 16'hC5D7, 16'hCE58, 16'hC618, 16'hC618, 16'hC618, 16'hC618, 16'hC618, 16'hC617, 16'hD699, 16'hACD3, 16'h4042, 16'hBD96, 16'hEF1C, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71D, 16'hC65A, 16'hC65A, 16'hC65A, 16'hEF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hB555, 16'h6A8A, 16'h6A4A, 16'h72CB, 16'hA492, 16'hC5D7, 16'hCE18, 16'hD69A, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hDE9B, 16'hA4D3, 16'h4083, 16'hBD96, 16'hCE59, 16'hC618, 16'hC618, 16'hCE18, 16'hCE18, 16'hD659, 16'hCDD7, 16'hACD3, 16'h9C10, 16'h9C51, 16'hA492, 16'hA492, 16'h4186, 16'h8B8E, 16'h4945, 16'h9451, 16'hB595, 16'h9CD2, 16'h000, 16'hA4D3, 16'hCE59, 16'hC618, 16'hC658, 16'hCE18, 16'hC618, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hC618, 16'hCE59, 16'hB555, 16'h5208, 16'hBD96, 16'hBDD7, 16'hB595, 16'h83CF, 16'h4145, 16'h83CE, 16'hBDD6, 16'h9C92, 16'h9C51, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hDE9A, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE59,
        16'hCE58, 16'hCE59, 16'hCE18, 16'hA4D2, 16'h59C7, 16'h830C, 16'hB515, 16'hD659, 16'hD659, 16'hCE59, 16'hCE59, 16'hCE19, 16'hCE19, 16'hCE18, 16'hCE18, 16'hCE18, 16'hCE18, 16'hCE59, 16'hBD96, 16'hA492, 16'hACD4, 16'hCE18, 16'hCE18, 16'hCE18, 16'hCE18, 16'hC618, 16'hC618, 16'hC617, 16'hCE58, 16'hB555, 16'h3843, 16'h2800, 16'h4985, 16'h6248, 16'h834D, 16'hB515, 16'hD659, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF9E, 16'hE75D, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hB4D4, 16'h6187, 16'h7B0C, 16'hD618, 16'hF6DC, 16'hC596, 16'hD658, 16'hDEDB, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD65A, 16'hD659, 16'hDE9A, 16'h9410, 16'h8B8E, 16'hCE59, 16'hC618, 16'hCE18, 16'hC618, 16'hC618, 16'hCE59, 16'hBD96, 16'h940F, 16'hA492, 16'hC597, 16'hCE18, 16'hCDD8, 16'hC5D7, 16'h628A, 16'h000,
        16'h9491, 16'hAD55, 16'hB595, 16'h9450, 16'h5A8A, 16'hC618, 16'hC658, 16'hCE58, 16'hCE58, 16'hCE18, 16'hCE18, 16'hCE58, 16'hC618, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE59, 16'hCE18, 16'h72CA, 16'h9491, 16'hBDD6, 16'hB595, 16'hBDD6, 16'hBDD7, 16'hB596, 16'h630B, 16'h840F, 16'hB596, 16'h7B0B, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hD69A, 16'hCE59, 16'hCE59, 16'hCE58, 16'hCE99, 16'hCE58, 16'h9C51, 16'h4904, 16'h834D, 16'hAC93, 16'hA452, 16'hA492, 16'hC596, 16'hD659, 16'hD659, 16'hCE19, 16'hCE19, 16'hCE19, 16'hCE18, 16'hCE59, 16'hCE18, 16'hCE18, 16'hCE19, 16'hBD56, 16'hA492, 16'hB555, 16'hCE18, 16'hC618, 16'hC618, 16'hC618, 16'hC618, 16'hC617, 16'hCE59, 16'h9411, 16'h8C0F, 16'hD659, 16'hBDD7, 16'hA4D3, 16'h83CF, 16'h7B4D, 16'h5A08, 16'h61C7, 16'h9410, 16'hCE18, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCDD7, 16'h69C8, 16'hA492, 16'hF71D, 16'hFF9E, 16'hEE9B, 16'hDE59, 16'hAC93, 16'hCE18, 16'hDE9A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hDE9A, 16'h838E, 16'h9410, 16'hCE59, 16'hC618, 16'hC618, 16'hC618, 16'hCE59, 16'hC5D7, 16'h9410, 16'hBD55, 16'hD619, 16'hD659, 16'hD659, 16'hCE18, 16'hD618, 16'h8B8E, 16'h62CB, 16'hB595, 16'hB595, 16'hB596, 16'h7B4C, 16'h9CD2, 16'hCE59, 16'hC618, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE18, 16'hCE58, 16'hC658, 16'hCE58, 16'hCE59, 16'hCE18, 16'hCE59, 16'hAD14, 16'h5A48, 16'hBDD6, 16'hB5D6, 16'hB5D6, 16'hBDD6, 16'hBDD6, 16'hBDD7, 16'hB596, 16'h5A89, 16'hAD13, 16'h838D, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hDE9A, 16'hCE59, 16'hCE59, 16'hCE18, 16'h8B4D, 16'h4883, 16'hBD15, 16'hD619, 16'hCDD7, 16'hC596, 16'hB4D4, 16'hA452, 16'hBD55, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hCE59, 16'hCE18, 16'hCE59, 16'hCE58, 16'hCE58, 16'hD619, 16'hB515, 16'hA492, 16'hBD96, 16'hCE18, 16'hC618, 16'hC618, 16'hC618, 16'hC618, 16'hC5D7, 16'h6208, 16'hAD14, 16'hDEDB, 16'hD69A, 16'hC5D8, 16'hB515, 16'hD69A, 16'hD659, 16'hB515, 16'h838F, 16'h5986, 16'h59C7, 16'hACD3, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h8B4E, 16'h830D, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hC596, 16'hC555, 16'hD618, 16'hB4D4, 16'hDE9A, 16'hDE9A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hDE9A, 16'h838E, 16'h9C11, 16'hD659, 16'hC618, 16'hCE18,
        16'hCE18, 16'hC5D7, 16'h9C51, 16'hBD55, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hCE18, 16'hDE59, 16'h9C11, 16'h49C7, 16'hB595, 16'hB596, 16'hBDD6, 16'h7B4C, 16'h9C91, 16'hCE59, 16'hC618, 16'hC618, 16'hCE18, 16'hCE18, 16'hCE58, 16'hCE58, 16'hC658, 16'hC658, 16'hCE58, 16'hCE59, 16'hCE19, 16'h72CB, 16'h9C91, 16'hC617, 16'hBDD7, 16'hBDD7, 16'hBDD7, 16'hC617, 16'hC617, 16'hC658, 16'h9451, 16'h7B8E, 16'h9451, 16'hAD14, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5E, 16'hDEDB, 16'hC596, 16'h5145, 16'h7ACC, 16'hD5D7, 16'hDE9A, 16'hD65A, 16'hDE9A, 16'hDE9A, 16'hD659, 16'hBD15, 16'hA452, 16'hBD55, 16'hD659, 16'hD659, 16'hD659, 16'hCE59, 16'hCE18, 16'hD659, 16'hCE59, 16'hCE18, 16'hCE59, 16'hCDD8, 16'hACD3, 16'hACD3, 16'hC5D7, 16'hCE18, 16'hC618, 16'hC618, 16'hCE59, 16'hA492, 16'h6A8A, 16'hD659, 16'hD69A,
        16'hD65A, 16'hBD55, 16'hA452, 16'hD659, 16'hCE18, 16'hCE18, 16'hDE9A, 16'hD659, 16'hAD13, 16'h6A8A, 16'h3000, 16'h9451, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE5A, 16'h7A09, 16'hBD15, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hABD0, 16'hE65A, 16'hD5D8, 16'hBD55, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hDE9A, 16'hDE9A, 16'h8B8E, 16'h9C51, 16'hD659, 16'hC618, 16'hCE18, 16'hCE18, 16'hA452, 16'hACD4, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hD619, 16'hD659, 16'hC596, 16'h5A08, 16'h62CB, 16'hB596, 16'hC618, 16'h8C0F, 16'h8C0F, 16'hCE59, 16'hC618, 16'hCE18, 16'hC618, 16'hCE18, 16'hCE18, 16'hCE59, 16'hCE58, 16'hCE58, 16'hC658, 16'hCE59, 16'hB555, 16'h5A07, 16'hC5D6, 16'hBDD7, 16'hBDD7, 16'hBDD7, 16'hC617, 16'hBDD6, 16'hAD55, 16'hCE18, 16'hAD54, 16'h7B8D, 16'hAD14, 16'h7B4D, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAC92, 16'h3800, 16'hA492, 16'hDE5A, 16'hDE9A, 16'hD65A, 16'hD65A, 16'hD65A, 16'hD659, 16'hDE9A, 16'hD659, 16'hB4D4, 16'hA452, 16'hBD56, 16'hD659, 16'hD659, 16'hD659, 16'hCE59, 16'hCE18, 16'hCE59, 16'hCE59, 16'hCE18, 16'hCE19, 16'hC596, 16'hA492, 16'hB555, 16'hCE18, 16'hC618, 16'hCE58, 16'hC5D7, 16'h59C7, 16'hAD14, 16'hDE9B, 16'hD659, 16'hD65A, 16'hB515, 16'hB555, 16'hD65A, 16'hAD14, 16'hB555, 16'hDE9A, 16'hD69A, 16'hDE9A, 16'hD659, 16'hB555, 16'h6249, 16'h2000, 16'hBD55, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC596, 16'h7A8B, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEE9B, 16'hCD56, 16'hFF1D, 16'hD5D8, 16'hCD97, 16'hDEDB,
        16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hD69A, 16'hDE9A, 16'h8BCF, 16'h9410, 16'hD659, 16'hCE18, 16'hCE19, 16'hB514, 16'hA452, 16'hCE19, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hDE5A, 16'hDE18, 16'hB412, 16'h3000, 16'h5A89, 16'hBDD7, 16'hAD54, 16'h6ACA, 16'hCE18, 16'hCE18, 16'hCE18, 16'hCE18, 16'hCE59, 16'hCE59, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE59, 16'hCE59, 16'h8B8E, 16'h83CF, 16'hC618, 16'hBDD7, 16'hBDD7, 16'hBE17, 16'hC617, 16'h7B8E, 16'h5A89, 16'hAD14, 16'hC5D7, 16'h734C, 16'hBD96, 16'h628A, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'h7A8A, 16'h830D, 16'hD619, 16'hEEDC, 16'hDE9A, 16'hDE5A, 16'hD65A, 16'hD65A, 16'hD659, 16'hD659, 16'hD659, 16'hDE9A, 16'hD619, 16'hAC93, 16'hA452, 16'hCDD8, 16'hD659, 16'hD659, 16'hD659, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE18,
        16'hCE18, 16'hD619, 16'hB555, 16'hACD3, 16'hC5D7, 16'hCE19, 16'hD659, 16'h93CF, 16'h72CB, 16'hDE9A, 16'hD69A, 16'hD69A, 16'hCE19, 16'h9C11, 16'hCDD8, 16'hD659, 16'hA492, 16'hC5D7, 16'hDE9A, 16'hD69A, 16'hD65A, 16'hD69A, 16'hDE9A, 16'hD69A, 16'hA4D3, 16'h3000, 16'h6208, 16'hCE17, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB4D4, 16'h938E, 16'hF75D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDDD8, 16'hEEDC, 16'hFFDF, 16'hE65A, 16'hE69B, 16'hE6DB, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hD69A, 16'hDE9A, 16'h9410, 16'h838E, 16'hD659, 16'hCE59, 16'hC596, 16'h93D0, 16'hC597, 16'hD659, 16'hD619, 16'hD659, 16'hD659, 16'hD659, 16'hDE9A, 16'hDE59, 16'hC514, 16'hAC11, 16'hC515, 16'hD598, 16'h8B8E, 16'h6248, 16'hBD96, 16'h730B, 16'hB555, 16'hCE59, 16'hCE18, 16'hCE18, 16'hCE18, 16'hCE58, 16'hCE58, 16'hCE18, 16'hCE58, 16'hCE59, 16'hC5D7, 16'h5A07, 16'hB595, 16'hC618, 16'hBDD7,
        16'hC617, 16'hC618, 16'hBDD6, 16'h734C, 16'hA4D3, 16'h83CF, 16'hBDD7, 16'h730C, 16'hC5D7, 16'h6ACB, 16'hCDD8, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hB4D3, 16'h82CC, 16'hCDD8, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'hF75D, 16'hEF1C, 16'hEF1C, 16'hEF1D, 16'hEF1C, 16'hE6DC, 16'hDE9A, 16'hD65A, 16'hDE9A, 16'hCDD8, 16'hAC52, 16'hBD14, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hCE59, 16'hCE18, 16'hCE18, 16'hCE18, 16'hCE59, 16'hC5D7, 16'hAD14, 16'hB555, 16'hD619, 16'hC596, 16'h6187, 16'hBD96, 16'hDE9B, 16'hD65A, 16'hDE9A, 16'hB515, 16'hAC93, 16'hDE9A, 16'hCE18, 16'hA492, 16'hD659, 16'hDE9A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD65A, 16'hD69A, 16'hDE9A, 16'hCE18, 16'h8C10, 16'h000, 16'h9C91, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA451, 16'hA410, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hCD56, 16'hF75E, 16'hFFDF, 16'hEEDC, 16'hF71D, 16'hE6DB, 16'hE6DB, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hD69A, 16'hDE9A, 16'hB4D4, 16'h6A09, 16'hCE18, 16'hD659, 16'hA492, 16'hB4D4, 16'hD65A, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hDE5A, 16'hB493, 16'hBD15, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB514, 16'h59C6, 16'h5A07, 16'h840F, 16'hC658, 16'hC618, 16'hCE58, 16'hCE58, 16'hCE18, 16'hCE58, 16'hCE58, 16'hCE58, 16'hD659, 16'hA491, 16'h6B0C, 16'hC618, 16'hC617, 16'hBE17, 16'hC618, 16'hC618, 16'hC618, 16'h840F, 16'h62CB, 16'h9C92, 16'hBDD7, 16'h734D, 16'hC617, 16'h940F, 16'hAC93, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hCDD7, 16'h830C, 16'hA410, 16'hE65A, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hF75E, 16'hEF1C, 16'hE6DB, 16'hC556, 16'hAC92, 16'hCDD7, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hCE18, 16'hCE18, 16'hCE58, 16'hCE18, 16'hC5D7, 16'hB555, 16'hCDD8, 16'h6A8A, 16'h9C11, 16'hDE9A, 16'hD69A, 16'hD69A, 16'hCE18, 16'hA452, 16'hCDD8, 16'hDE9A, 16'hBD55, 16'hACD4, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hDE9A, 16'hBD96, 16'h6209, 16'h6A49, 16'hE6DC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9BD0, 16'hAC93, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'hD597, 16'hFFDF, 16'hFF9F, 16'hEE9B, 16'hFF9E, 16'hF71D, 16'hE6DB, 16'hE6DB, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hC596, 16'h6187, 16'hBD96, 16'hC5D7, 16'h9C51, 16'hCE18, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hDE5A, 16'hBCD4, 16'hC556, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCDD7, 16'h5001, 16'h6249, 16'hCE18, 16'hCE59,
        16'hCE18, 16'hCE58, 16'hCE18, 16'hCE59, 16'hCE59, 16'hCE59, 16'hD618, 16'h6A8A, 16'hAD14, 16'hCE59, 16'hC617, 16'hC618, 16'hC618, 16'hBDD7, 16'hCE58, 16'hBDD7, 16'hAD54, 16'hC658, 16'hBDD7, 16'h7B8E, 16'hC5D7, 16'hB514, 16'h7ACB, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hCD97, 16'h7208, 16'h830C, 16'hE6DB, 16'hFF9E, 16'hD5D8, 16'hCD56, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF79E, 16'hE69B, 16'hAC93, 16'hB4D4, 16'hD659, 16'hD659, 16'hD659, 16'hCE59, 16'hCE18, 16'hCE18, 16'hCE18, 16'hCE18, 16'hCE19, 16'hCE18, 16'hD619, 16'hA452, 16'h6249, 16'hD659, 16'hDE9A, 16'hD69A, 16'hDE5A, 16'hAC93, 16'hB515, 16'hDE9A, 16'hD659, 16'hAC93, 16'hC5D7, 16'hDEDB, 16'hDE9A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hDE9A, 16'hD659, 16'h838E, 16'h4801, 16'hD65A,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA410, 16'hB493, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE61A, 16'hE65A, 16'hFFDF, 16'hFF9F, 16'hE65A, 16'hFF9F, 16'hFFDF, 16'hEEDC, 16'hE6DB, 16'hDEDB, 16'hDE9A, 16'hDE9A, 16'hDE9B, 16'hD659, 16'hCDD7, 16'h834D, 16'hA451, 16'hAC92, 16'hB514, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hDE9A, 16'hCD96, 16'hBCD4, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE5A, 16'h7209, 16'h7B0C, 16'hC5D7, 16'hD659, 16'hC618, 16'hCE18, 16'hCE58, 16'hCE58, 16'hD699, 16'hBD55, 16'h628A, 16'hC618, 16'hC658, 16'hC618, 16'hC617, 16'hCE59, 16'hEF1C, 16'hF79E, 16'hEF5D, 16'hCE99, 16'hC658, 16'hC617, 16'h83CE, 16'hBDD6, 16'hC5D7, 16'h724A, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hCD97, 16'h824A, 16'h7A09, 16'hD5D8, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hF75D, 16'hD597, 16'hD557, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hC596, 16'hA452, 16'hCDD7, 16'hD699, 16'hD659, 16'hD659, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE18, 16'hCE18, 16'hCE59, 16'hC5D7, 16'h5003, 16'hBD96, 16'hDEDB, 16'hD69A, 16'hDE9A, 16'hC596, 16'hA452, 16'hD659, 16'hDE9A, 16'hC556, 16'hAC93, 16'hDE9A, 16'hDE9A, 16'hD69A, 16'hD69A, 16'hDE9A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'h9C91, 16'h3800, 16'hCDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD15, 16'hA410, 16'hFFDF, 16'hF75D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD598, 16'hEE9B, 16'hFFDF, 16'hFF9E, 16'hE65A, 16'hFF9F, 16'hFFDF, 16'hF79E, 16'hE6DB, 16'hE6DB, 16'hDEDB, 16'hDE9A, 16'hE6DB, 16'hCE18, 16'hC597, 16'hA493, 16'h5986, 16'h9C10, 16'hCE18, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hDE5A, 16'hD619, 16'hB493, 16'hEEDC,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hEEDC, 16'hD597, 16'h7A8B, 16'h5003, 16'hB514, 16'hE69A, 16'hD65A, 16'hCE18, 16'hCE18, 16'hD659, 16'h8B8E, 16'h8C10, 16'hCE59, 16'hC618, 16'hC618, 16'hDE9B, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hDEDB, 16'hC617, 16'h7BCE, 16'hBDD6, 16'hCE18, 16'h7ACB, 16'hCD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'hBD14, 16'h7A4A, 16'h7A8A, 16'hD5D7, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hCD56, 16'hDDD8, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'hAC93, 16'hB515, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hCE59, 16'hCE18, 16'hCE18, 16'hD659, 16'h830C, 16'h93CF, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hD618, 16'hA452, 16'hCDD8, 16'hDE9B, 16'hD619, 16'hAC93, 16'hCDD8, 16'hDEDB, 16'hDE9A, 16'hDE9A, 16'hDE9A,
        16'hDE9A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hDE9A, 16'hA492, 16'h2800, 16'hC597, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCDD7, 16'h9B8E, 16'hFF9E, 16'hF71D, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hD597, 16'hF71D, 16'hFFDF, 16'hFF9E, 16'hE69A, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hEF1D, 16'hE6DB, 16'hE6DB, 16'hDE9A, 16'hE6DB, 16'hC596, 16'hCDD8, 16'hCE18, 16'h4800, 16'hA452, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hD65A, 16'hDE9A, 16'hBCD4, 16'hCD97, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hDE19, 16'hEEDB, 16'hFFDF, 16'hFF9F, 16'hC596, 16'h7208, 16'hA3CF, 16'hE69A, 16'hF75D, 16'hE71C, 16'hCDD8, 16'h59C6, 16'hB595, 16'hCE18, 16'hC618, 16'hDE9B, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h7B8E, 16'hBDD6, 16'hC618, 16'h9C51, 16'hAC11, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hDE59,
        16'hB514, 16'h930C, 16'h6884, 16'h930D, 16'hCD56, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69B, 16'hC4D5, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hCD97, 16'hA492, 16'hCDD8, 16'hD659, 16'hD659, 16'hD659, 16'hCE19, 16'hCE18, 16'hCE18, 16'hD659, 16'h9C10, 16'h7B0C, 16'hD659, 16'hDE9B, 16'hD69A, 16'hDE5A, 16'hB4D4, 16'hBD56, 16'hE69B, 16'hDE9A, 16'hBD55, 16'hBD56, 16'hDEDB, 16'hDEDA, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hDE9A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'h9C51, 16'h2800, 16'hCDD8, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD618, 16'h8B0C, 16'hFF5E, 16'hF75D, 16'hDE19, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hD557, 16'hFF5E, 16'hFFDF, 16'hFF5E, 16'hEE9B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hE71C, 16'hE6DB, 16'hE6DB, 16'hE6DB, 16'hC556, 16'hCE18,
        16'hE69B, 16'h8B4E, 16'h93CF, 16'hDE5A, 16'hD659, 16'hD659, 16'hD659, 16'hDE9A, 16'hD618, 16'hBC94, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hDE19, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hB4D3, 16'h7249, 16'h9C10, 16'hE69A, 16'hCD56, 16'h7B8E, 16'hD659, 16'hC618, 16'hD69A, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DC, 16'h83CF, 16'hCE18, 16'hD659, 16'hCE17, 16'h7A09, 16'hEF1C, 16'hFF9E, 16'hEE9B, 16'hCD97, 16'hBC93, 16'h9B4E, 16'h928B, 16'hA38E, 16'hB4D3, 16'hD618, 16'hF71D, 16'hFF5E, 16'hDDD8, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hCD97, 16'hCD57, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hEF1C, 16'hD618, 16'hAC92, 16'hBD55, 16'hD659, 16'hD659, 16'hD659, 16'hCE19, 16'hCE18, 16'hDE59, 16'h9C10, 16'h59C7, 16'hD618, 16'hDE9B, 16'hDE9A, 16'hDE9A,
        16'hBD56, 16'hB4D4, 16'hDE9A, 16'hE69B, 16'hCDD7, 16'hB514, 16'hDE9A, 16'hDEDB, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hCE58, 16'hACD3, 16'h8B4E, 16'h4000, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h7186, 16'hEEDC, 16'hFFDF, 16'hDE19, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD597, 16'hFF5E, 16'hFFDF, 16'hF71D, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hE6DC, 16'hE6DB, 16'hDE9A, 16'hC555, 16'hD659, 16'hDE9B, 16'hAC92, 16'h6185, 16'hC597, 16'hD659, 16'hD659, 16'hD659, 16'hDE9A, 16'hC515, 16'hD5D8, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9B, 16'hDDD8, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69B, 16'hA411, 16'h828B, 16'h6145, 16'h72CB, 16'hA492, 16'hAD14, 16'hE6DB, 16'hF71D, 16'hE69B, 16'hCD97, 16'hAC92, 16'h9C11, 16'hA451, 16'hBD14, 16'hD5D8, 16'hBD55, 16'h6A49,
        16'h9C10, 16'h8B4D, 16'h7289, 16'h000, 16'h71C8, 16'h92CC, 16'h92CC, 16'hA38F, 16'hC515, 16'hDE59, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65A, 16'hDD97, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'hC4D5, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hE6DB, 16'hDE5A, 16'hDE9A, 16'hBD15, 16'hACD3, 16'hCE18, 16'hD659, 16'hD659, 16'hCE59, 16'hD659, 16'hA451, 16'h61C8, 16'hCDD7, 16'hE6DB, 16'hDE9A, 16'hE69B, 16'hD619, 16'hAC52, 16'hD659, 16'hE6DB, 16'hD659, 16'hBD15, 16'hDE9A, 16'hE71C, 16'hE6DB, 16'hDEDB, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hD69A, 16'hD69A, 16'hDE9A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hDE9A, 16'hD69A, 16'hD69A, 16'hDE9A, 16'hD659, 16'hA493, 16'hACD3, 16'hCE18, 16'h8B8F, 16'h59C7, 16'hEF5C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'h828B, 16'hDE5A, 16'hFFDF, 16'hF75E, 16'hE65A, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hDDD9, 16'hF75D, 16'hFFDF,
        16'hF71E, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1D, 16'hE6DC, 16'hE69A, 16'hCD96, 16'hDE5A, 16'hDE9A, 16'hC596, 16'h830C, 16'h8B8E, 16'hDE59, 16'hCE59, 16'hD65A, 16'hD5D8, 16'hBCD4, 16'hEF1D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hDDD8, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1D, 16'hFF5E, 16'hFFDF, 16'hFF5E, 16'hE69B, 16'hBD14, 16'h9BCF, 16'h938E, 16'h7209, 16'h7A09, 16'h8B0D, 16'h934D, 16'hB4D3, 16'hCDD8, 16'hCDD7, 16'hB493, 16'h9B8F, 16'h8B4D, 16'h938F, 16'hA452, 16'hACD3, 16'hC556, 16'hCDD7, 16'hDE5A, 16'hEF1C, 16'hF71D, 16'hDDD8, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hD556, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hCD57, 16'hD5D8, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hEF1D, 16'hDE9A, 16'hDE5A, 16'hDE5A, 16'hDE9A, 16'hCDD7, 16'hACD3,
        16'hC5D7, 16'hD659, 16'hD659, 16'hDE59, 16'hA451, 16'h61C6, 16'hCDD7, 16'hE6DB, 16'hDE9A, 16'hDE9B, 16'hE6DB, 16'hC556, 16'hCD97, 16'hEF5D, 16'hF75D, 16'hEEDC, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hF75E, 16'hF75D, 16'hEF1D, 16'hE71C, 16'hDEDB, 16'hDE9A, 16'hD69A, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hACD4, 16'hAD14, 16'hD65A, 16'hCE18, 16'hA492, 16'h6A49, 16'h93D0, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA411, 16'hC555, 16'hFFDF, 16'hDE19, 16'hF71D, 16'hEEDC, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9C, 16'hF75D, 16'hFFDF, 16'hF6DC, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hEF1C, 16'hE69B, 16'hD5D7, 16'hDE9A, 16'hD65A, 16'hD5D8, 16'hCD97, 16'h61C6, 16'hC596, 16'hD65A, 16'hDE9A, 16'hC555, 16'hCD97, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'hDDD8, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hEE9B, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hEE9B, 16'hC515, 16'hF71C, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9B, 16'hEE9B, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hD597, 16'hE65A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE19, 16'hE619, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE19, 16'hC4D5, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hEEDC, 16'hDE9A, 16'hDE5A, 16'hDE9A, 16'hDE5A, 16'hDE9A, 16'hCE18, 16'hACD3, 16'hBD96, 16'hD65A, 16'hD619, 16'hA451, 16'h724A, 16'hCE17, 16'hE6DB, 16'hDE9A, 16'hE6DB, 16'hE6DB, 16'hEF1C, 16'hF71D, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hF75D, 16'hE71C, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hDEDA, 16'hDE9A, 16'hBD55, 16'hA492, 16'hD659, 16'hDE9A, 16'hACD3, 16'h9C92, 16'hC5D7, 16'h5947, 16'hC596, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD618, 16'h938E, 16'hFFDF, 16'hF71C, 16'hCD56, 16'hFF9E, 16'hEE9B,
        16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hFF5E, 16'hFF9F, 16'hE65A, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hEEDC, 16'hE69B, 16'hE6DC, 16'hD659, 16'hCDD7, 16'hE6DB, 16'h9BD0, 16'h7ACC, 16'hD659, 16'hDE5A, 16'hBCD4, 16'hE65A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hDDD8, 16'hEE9B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hEE9B, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD57, 16'hDE5A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hCD56, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hDDD8, 16'hE619, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9B, 16'hD557, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'hC4D5, 16'hEEDC, 16'hFFDF,
        16'hFFDF, 16'hFF9F, 16'hF75E, 16'hE6DB, 16'hDE5A, 16'hDE5A, 16'hDE5A, 16'hDE5A, 16'hDE59, 16'hDE5A, 16'hD659, 16'hBD55, 16'hC596, 16'hCDD8, 16'h8B8E, 16'h6A49, 16'hD5D8, 16'hE6DB, 16'hE6DB, 16'hE6DC, 16'hF75D, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hE71C, 16'hDEDB, 16'hDEDB, 16'hCE18, 16'hACD3, 16'hCE18, 16'hD65A, 16'hB515, 16'h9C10, 16'hC617, 16'hDEDB, 16'hA492, 16'h50C4, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h82CB, 16'hF75D, 16'hFFDF, 16'hCD56, 16'hE65A, 16'hFFDF, 16'hE65A, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF1D, 16'hF71D, 16'hFF9E, 16'hEE9B, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hE69B, 16'hF75D, 16'hF75E, 16'hD618, 16'hD618, 16'hE6DC, 16'hD5D8, 16'h6187, 16'hB514, 16'hDE59, 16'hB4D4, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hD557, 16'hFF5E, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hEE9B, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hC4D4, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hD557, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE619, 16'hDDD8, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF6DD, 16'hCD16, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hCD16, 16'hDE19, 16'hFFDF, 16'hFF9F, 16'hF75E, 16'hE6DB, 16'hDE9A, 16'hDE9A, 16'hDE5A, 16'hDE5A, 16'hDE5A, 16'hDE5A, 16'hD659, 16'hD65A, 16'hD619, 16'hBD15, 16'h6A08, 16'h830C, 16'hD619, 16'hEF1D, 16'hF75D, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hE61A, 16'hFF5E, 16'hFF9F, 16'hEEDC, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hE6DB,
        16'hCDD8, 16'hCE18, 16'hDE9B, 16'hC597, 16'h9410, 16'hC597, 16'hDE9A, 16'hD6DA, 16'hCE59, 16'h61C8, 16'hAC92, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h93CF, 16'hD619, 16'hFFDF, 16'hFFDF, 16'hD5D8, 16'hE69A, 16'hFFDF, 16'hE65A, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9C, 16'hEE9B, 16'hFF9F, 16'hF6DC, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65A, 16'hF75D, 16'hFFDF, 16'hE69A, 16'hDE9A, 16'hE6DC, 16'hE6DC, 16'hB514, 16'h5986, 16'hBD14, 16'hC556, 16'hFF5E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65A, 16'hDDD9, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9B, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69B, 16'hCD56, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'hDDD9, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE5A, 16'hDD98, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hCD56, 16'hEE9B,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD5D8, 16'hCD57, 16'hFF5E, 16'hF75D, 16'hE69B, 16'hDE5A, 16'hDE5A, 16'hDE5A, 16'hDE5A, 16'hDE5A, 16'hDE5A, 16'hDE59, 16'hDE9A, 16'hDE5A, 16'hA452, 16'h71C8, 16'hB4D4, 16'hF75D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65A, 16'hE61A, 16'hFFDF, 16'hF6DC, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69B, 16'hD5D8, 16'hEF1C, 16'hE6DB, 16'hD619, 16'hA452, 16'hBD96, 16'hDEDA, 16'hD69A, 16'hD69A, 16'hDEDA, 16'hACD4, 16'h4800, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCDD7, 16'h9BCF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDDD8, 16'hE65A, 16'hFFDF, 16'hE65A, 16'hEE9B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDDD8, 16'hEE9B, 16'hFF9F, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hD597, 16'hF75D, 16'hFFDF, 16'hFF5E, 16'hF75E, 16'hE71C, 16'hE6DB, 16'hE69B, 16'h9C10, 16'h7A8A, 16'hBD15,
        16'hEEDC, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hD597, 16'hEE9B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hE65A, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE19, 16'hDDD8, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9B, 16'hDE19, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9B, 16'hDD97, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hD5D8, 16'hDDD8, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65A, 16'hC515, 16'hDE5A, 16'hDE9B, 16'hDE5A, 16'hDE9A, 16'hDE5A, 16'hDE5A, 16'hDE59, 16'hDE59, 16'hDE5A, 16'hDE9A, 16'hCDD7, 16'h8B4D, 16'h830C, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF6DD, 16'hDDD8, 16'hFF9F, 16'hFF5E, 16'hEE9B, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65B, 16'hC516, 16'hF71D, 16'hFFDF, 16'hF75D, 16'hB514, 16'hB555, 16'hDEDB, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD659, 16'h728A, 16'h9C51, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'h828A, 16'hEF1C, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDDD9, 16'hE619, 16'hFFDF, 16'hEE9B, 16'hE65A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hCD56, 16'hF75D, 16'hFF9F, 16'hF6DC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hD5D7, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hE6DC, 16'hE6DC, 16'hDE5A, 16'h7A8A, 16'h82CC, 16'hDE19, 16'hF71D, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF71D, 16'hD557, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9C, 16'hE69B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hD557, 16'hE69B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69A, 16'hE619, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDC,
        16'hD557, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65A, 16'hCD16, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hB493, 16'hC597, 16'hDE9A, 16'hDE9A, 16'hDE5A, 16'hDE5A, 16'hDE5A, 16'hD659, 16'hDE5A, 16'hDE5A, 16'hA452, 16'h6906, 16'hB4D3, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hDD98, 16'hF71D, 16'hFFDF, 16'hF71D, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDB, 16'hCD16, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hC555, 16'hD69A, 16'hDEDA, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD699, 16'hDE9A, 16'hB514, 16'h3000, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9B90, 16'hC556, 16'hFF5E, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hE65A, 16'hE619, 16'hFFDF, 16'hE69B, 16'hE65A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9B, 16'hCD56, 16'hFFDF, 16'hFF9F, 16'hFF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hF71D, 16'hEE5B, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hDEDB, 16'hE6DC, 16'hD618, 16'h5946, 16'hA451, 16'hE69A, 16'hF71D, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE65B, 16'hD597, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hE619, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hC4D5, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65A, 16'hDE19, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'hD557, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1D, 16'hCCD5, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hE69B, 16'hB494, 16'hC556, 16'hDE9A, 16'hDE5A, 16'hDE9A, 16'hDE5A, 16'hDE5A, 16'hDE9A, 16'hC556, 16'h828B, 16'h830C, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hE65A, 16'hE65A, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF6DC, 16'hD597, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hE65A, 16'hEEDC, 16'hE71C, 16'hDE9A, 16'hDE9A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD659, 16'h6A8A, 16'hACD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD618, 16'h8B0D, 16'hF71D, 16'hCD16, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hE65A, 16'hDE19, 16'hFFDF, 16'hE69B, 16'hEE9B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDDD8, 16'hD597, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hF6DD, 16'hFFDF, 16'hEE9B, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1D, 16'hDEDB, 16'hE6DC, 16'hBD15, 16'h5082, 16'hBCD4, 16'hE69B, 16'hEF1D, 16'hFF9F, 16'hFF9F, 16'hDE19, 16'hDDD9, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5D, 16'hDDD8, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'hCCD5, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65A,
        16'hDE5A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hD557, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hCD16, 16'hDE19, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hE6DB, 16'hDE5A, 16'hBD15, 16'hBD15, 16'hDE5A, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hD619, 16'hB492, 16'h7248, 16'h9BD0, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hDDD9, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hD598, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9B, 16'hE65A, 16'hFFDF, 16'hF75D, 16'hDE9B, 16'hDE9A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hDE9B, 16'hA4D3, 16'h59C7, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h828B, 16'hE65A, 16'hF71D, 16'hCD16, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hEE9B, 16'hDDD8, 16'hFFDF, 16'hDE19, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hD597, 16'hD5D7, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hFF9F, 16'hFFDF, 16'hE619, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hE6DC, 16'hDEDB, 16'hE6DB, 16'hB4D4, 16'h58C5, 16'hC555, 16'hE69B, 16'hEF1C, 16'hF75D, 16'hCD97, 16'hE65A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF6DC, 16'hDE19, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9B, 16'hCD16, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hDE19, 16'hE65A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hCD56, 16'hE65A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD598, 16'hD597, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF71D, 16'hE69A, 16'hDE59, 16'hDE5A, 16'hC555, 16'hBD15, 16'hDE5A, 16'hDE9A, 16'hDE59, 16'hC555, 16'h934D, 16'h8ACB, 16'hCDD7, 16'hF79E,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'hF71C, 16'hFFDF, 16'hF71D, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65B, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9B, 16'hDDD8, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hE6DB, 16'hDE9A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD619, 16'h61C7, 16'hCDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC556, 16'h9BCF, 16'hFFDF, 16'hFF9E, 16'hD598, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'hD597, 16'hFF5E, 16'hE65A, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hC4D4, 16'hDE19, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hE61A, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hDEDB, 16'hDEDB, 16'hE69B, 16'hB493, 16'h4000, 16'hB4D3, 16'hE6DC, 16'hDE9A, 16'hB493, 16'hE61A, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65A, 16'hDE19, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hE619, 16'hD557, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hDE19, 16'hDE19, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hD557, 16'hDE19, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65A, 16'hCCD5, 16'hF71D, 16'hFFDF, 16'hFF9E, 16'hF71D, 16'hE69B, 16'hDE5A, 16'hDE5A, 16'hDE9A, 16'hDE9A, 16'hCDD7, 16'hC556, 16'hDE19, 16'hC596, 16'hA410, 16'hB411, 16'hA34F, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hFFDF, 16'hFF5E, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65A, 16'hD557, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hDE9A, 16'hD69A, 16'hD69A,
        16'hD69A, 16'hD69A, 16'hD69A, 16'hDEDA, 16'h9C51, 16'h7B4D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h7188, 16'hDE59, 16'hFFDF, 16'hFF9F, 16'hCD97, 16'hEEDC, 16'hFFDF, 16'hFFDF,
        16'hF71D, 16'hD597, 16'hF71D, 16'hE69A, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hBC52, 16'hE69B, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hEE9C, 16'hFF9F, 16'hFF9F, 16'hEE5A, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1D, 16'hDE9B, 16'hE6DB, 16'hE6DB, 16'hBD15, 16'h6146, 16'hACD3, 16'hD618, 16'hBD15, 16'hDE19, 16'hF75D, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hD5D8, 16'hE65A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDD98, 16'hDD98, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE19, 16'hDDD8, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hD598, 16'hDDD9, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF6DD, 16'hCD15, 16'hE65A, 16'hEF1D, 16'hE69A, 16'hDE5A, 16'hDE5A, 16'hE65A, 16'hDE5A,
        16'hDE59, 16'hD5D8, 16'hC555, 16'hBCD3, 16'hAC51, 16'hB4D3, 16'hDDD8, 16'hD557, 16'hC494, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hE69A, 16'hFFDF, 16'hF71D, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hDDD8, 16'hD556, 16'hFF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hDEDB, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hDE9A, 16'hBD96, 16'h4903, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB4D4, 16'h9BD0, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hDE19, 16'hE69A, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hCD56, 16'hEE9B, 16'hEEDB, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hBC93, 16'hEEDB, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hE619, 16'hFF9F, 16'hFFDF, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hE6DC, 16'hE6DB, 16'hE6DB, 16'hEEDC, 16'hBD15, 16'h5040, 16'h938E, 16'hCD56, 16'hDE19,
        16'hDE9A, 16'hEEDC, 16'hF71D, 16'hFF9F, 16'hFF5E, 16'hCD56, 16'hEE9B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hD557, 16'hDDD9, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE659, 16'hD5D8, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hDDD9, 16'hD597, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hC515, 16'hBD15, 16'hD619, 16'hDE5A, 16'hDE5A, 16'hDE5A, 16'hD5D7, 16'hBD15, 16'hBCD4, 16'hAC51, 16'hC515, 16'hCD56, 16'hDDD8, 16'hE65B, 16'hEEDB, 16'hD597, 16'hE619, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD556, 16'hEE9B, 16'hFFDF, 16'hF6DC, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hE65A, 16'hFF5E, 16'hFFDF, 16'hFFDF,
        16'hEE9B, 16'hE65A, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD69A, 16'hD659, 16'h6208, 16'hB555, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hF75E, 16'h69C8, 16'hE69B, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'hEEDC, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hDDD8, 16'hEE9B, 16'hF71D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hEEDB, 16'hBC52, 16'hF71C, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hDDD8, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hE6DB, 16'hE6DC, 16'hD659, 16'hD618, 16'hD618, 16'h82CB, 16'h69C6, 16'hA451, 16'hD5D8, 16'hDE19, 16'hDE5A, 16'hEEDB, 16'hEE9B, 16'hC515, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hD516, 16'hDDD9, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65A, 16'hCD97, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE65A, 16'hCD16, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFF9F, 16'hF75D, 16'hE69B, 16'hC515, 16'hB4D4, 16'hDE59, 16'hE65A, 16'hCD57, 16'hAC52, 16'hAC52, 16'hC515, 16'hD5D7, 16'hD618, 16'hE69B, 16'hE69B, 16'hEEDB, 16'hEEDC, 16'hF71D, 16'hE619, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE619, 16'hD597, 16'hFFDF, 16'hF71D, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE19, 16'hE65A, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hD69A, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hCE19, 16'hCE18, 16'hDE9A, 16'h9410, 16'h730B, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD97, 16'h828A, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9B, 16'hC515, 16'hF71D, 16'hEE9B, 16'hE65A, 16'hF71D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hE69A, 16'hBC93, 16'hF71D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hD597, 16'hFF9F, 16'hF71D, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hE6DC, 16'hC597, 16'hD619, 16'hE6DC, 16'hD618, 16'hB493, 16'h7208, 16'h6A09, 16'hAC52, 16'hD5D7, 16'hE65A, 16'hD618, 16'hB493, 16'hE65A, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hCD16, 16'hDDD9, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9B, 16'hC516, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9B, 16'hC4D5, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF75D, 16'hEEDC, 16'hDE9B, 16'hE6DB, 16'hDE59, 16'hC515, 16'hC515, 16'hB452, 16'hA38F, 16'hB493, 16'hD5D8, 16'hE61A, 16'hE65A, 16'hEF1D, 16'hEEDC, 16'hEF1C, 16'hF75D, 16'hFFDF, 16'hF6DC, 16'hEE5A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hCD16, 16'hF71D, 16'hFFDF, 16'hEE9B, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF6DC, 16'hE619, 16'hFF9F, 16'hFFDF, 16'hF71D, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hDE9B, 16'hDE9A, 16'hD619, 16'hBD55, 16'hACD4, 16'hCE18, 16'hDE9B, 16'hB556, 16'h4040, 16'hE6DC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'h7ACB, 16'hB4D4, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'hF71C, 16'hB412, 16'hCD56, 16'hFF9F, 16'hEEDC, 16'hDE19, 16'hEEDC, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hE65A, 16'hBC93, 16'hF75D, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hD597, 16'hFF9F, 16'hE65A, 16'hEE9B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1D, 16'hC556, 16'hEEDC, 16'hF75D, 16'hDE9A, 16'hDE5A, 16'hDE19, 16'hB493, 16'h7A8A, 16'h8B0D, 16'hB4D4, 16'hC556, 16'hBC93, 16'hD5D8, 16'hE69A, 16'hE6DC, 16'hEF1C, 16'hF75D, 16'hFF9E, 16'hFF9F, 16'hFF9E, 16'hCD16, 16'hDDD8, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9C, 16'hC4D5, 16'hEEDC, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hEEDC, 16'hC4D5, 16'hDE19, 16'hFF9E, 16'hF75D, 16'hF75D, 16'hEF1D, 16'hEEDC, 16'hEF1C, 16'hEEDB, 16'hE65A, 16'hD5D8, 16'hBCD4, 16'h8A8C, 16'hA38F, 16'hCD56, 16'hD597, 16'hCD56, 16'hEEDC, 16'hD5D8, 16'hD5D8, 16'hEF1D, 16'hF75D, 16'hFF9F, 16'hFFDF, 16'hFF5E, 16'hDDD9, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE61A, 16'hDDD9, 16'hFFDF, 16'hF71C, 16'hE65A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hE65A, 16'hF71D, 16'hFFDF, 16'hFF9E, 16'hDE19, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hE6DB, 16'hCDD8, 16'hA492, 16'hA452, 16'hCDD7, 16'hDE9A, 16'hCE19, 16'hAD14, 16'h3000, 16'hCDD8, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69B, 16'h71C8, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE19, 16'hD598, 16'hE65A, 16'hA38F, 16'hF71C, 16'hFFDF, 16'hF71D, 16'hC516, 16'hE65A, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hEF1D, 16'hDE5A, 16'hC4D4, 16'hF75D, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hDDD8, 16'hFF9F, 16'hDE19, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hC556, 16'hF71D, 16'hFFDF, 16'hFF9E, 16'hE6DB, 16'hDE9A, 16'hDE19, 16'hD597, 16'hBCD4, 16'h7A4A, 16'h6A09, 16'h7209, 16'hB492, 16'hE659, 16'hE69B, 16'hE69B, 16'hDE9A, 16'hDE9A, 16'hE69B, 16'hE69B, 16'hC515, 16'hC515, 16'hE6DB, 16'hEEDC, 16'hEF1C, 16'hEF1C, 16'hEF1C, 16'hEEDC, 16'hEF1C, 16'hE69A, 16'hC515, 16'hD5D8, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDB, 16'hEEDB, 16'hE6DB, 16'hE69B, 16'hE69B, 16'hDE5A, 16'hC515, 16'hCD56, 16'hE6DB, 16'hEF1C, 16'hEF1C, 16'hEEDB, 16'hE659, 16'hCD97, 16'hAC92, 16'h9B4E, 16'h9B0E, 16'hBCD4, 16'hDE19, 16'hF71C, 16'hEE9B, 16'hAC51, 16'hCD97, 16'hF6DC, 16'hB493, 16'hDE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hDD98, 16'hF6DC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E,
        16'hD598, 16'hFF5E, 16'hFFDF, 16'hDE19, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hD597, 16'hDE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hDE19, 16'hBD14, 16'hC556, 16'hDE5A, 16'hDE9A, 16'hBD56, 16'h93D0, 16'hACD3, 16'h6ACB, 16'h9450, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAC92, 16'h9BD0, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF71D, 16'hDE18, 16'hFF5E, 16'hFF5E, 16'hB412, 16'hEEDC, 16'hFFDF, 16'hFF9F, 16'hDE19, 16'hE69A, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hEF1C, 16'hDE19, 16'hC515, 16'hF75D, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hEE9B, 16'hFF9F, 16'hEF1C, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD56, 16'hE65B, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF6DC, 16'hBD15, 16'hBD15, 16'hE69B, 16'hD598, 16'hB493, 16'hA411, 16'h828A, 16'h930C, 16'hAC92, 16'hCDD7, 16'hE65A, 16'hE69B, 16'hE69B, 16'hE69B, 16'hCD97, 16'hB4D3, 16'hDE59, 16'hDE9A, 16'hDE9A, 16'hDE9A,
        16'hDE9A, 16'hDE9A, 16'hE69A, 16'hE69A, 16'hC555, 16'hC556, 16'hE69A, 16'hE69A, 16'hDE9A, 16'hDE5A, 16'hDE5A, 16'hDE5A, 16'hDE5A, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hE69B, 16'hD5D8, 16'hCD56, 16'hE65A, 16'hD5D8, 16'hBCD4, 16'hA38F, 16'h9ACD, 16'h92CC, 16'hB453, 16'hDE19, 16'hFF5E, 16'hFFDF, 16'hFF9E, 16'hE69B, 16'hC555, 16'hB492, 16'hEE9C, 16'hE69B, 16'hBCD4, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hDDD8, 16'hEE9B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9B, 16'hE65A, 16'hFFDF, 16'hF71D, 16'hDDD9, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hB453, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hCD97, 16'hE69A, 16'hE69B, 16'hDE9A, 16'hD618, 16'hA493, 16'h9C51, 16'hC596, 16'hD69A, 16'h9C92, 16'h5A08,
        16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'h5043, 16'hC556, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hEE9B, 16'hFF5D, 16'hFFDF, 16'hFF9F, 16'hC4D4, 16'hDE5A, 16'hFFDF, 16'hFF9F, 16'hEEDC, 16'hE69B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hF75E, 16'hEEDC, 16'hDE19, 16'hCD55, 16'hF75D, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'hF75E, 16'hFFDF, 16'hFF5E, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD557, 16'hC515, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCD97, 16'hC555, 16'hD5D8, 16'hDE19, 16'hB4D4, 16'hC556, 16'hE659, 16'hC556, 16'h938E, 16'h7208, 16'h8B0D, 16'hAC51, 16'hC556, 16'hDE19, 16'hDE1A, 16'hCD56, 16'hDE59, 16'hE6DB, 16'hE6DB, 16'hE69A, 16'hE69B, 16'hE69A, 16'hDE9A, 16'hE69A, 16'hCDD8, 16'hBD55, 16'hDE5A, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE69B, 16'hE69B, 16'hE69B, 16'hDE59, 16'hD618, 16'hC556, 16'hB451, 16'h930D, 16'h934D, 16'h934E, 16'hB493, 16'hCD56, 16'hE69B, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hDE59, 16'hD5D8, 16'hCD56, 16'hDE19, 16'hFF9F, 16'hEEDB, 16'hDD97, 16'hFF9F, 16'hFFDF, 16'hF71D, 16'hDDD8, 16'hF6DC, 16'hFF5E, 16'hF71C, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9B, 16'hF75E, 16'hFFDF, 16'hEE9B, 16'hE65A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hE65B, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hF71D, 16'hFF9F, 16'hEF1D, 16'hBD55, 16'hA492, 16'hBD96, 16'hD69A, 16'hD69A, 16'hDEDA, 16'hBD96, 16'h3800, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69B, 16'h9C11, 16'h6188, 16'hEEDC, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hF71C, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hCD97, 16'hD5D8, 16'hF75D, 16'hF71D, 16'hE65A, 16'hC4D5, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1D, 16'hE6DC, 16'hD618, 16'hCD56, 16'hF75D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hEEDB, 16'hFF9F, 16'hFFDF, 16'hF71D, 16'hD597, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hE65A, 16'hEE9B, 16'hC4D5, 16'hF71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEE9C, 16'hF6DC, 16'hCD97, 16'hEE9B, 16'hD5D8, 16'hB493, 16'hBD55, 16'hF6DC,
        16'hFF5E, 16'hE69B, 16'hC556, 16'h938F, 16'h828B, 16'h828B, 16'h9B4F, 16'hAC12, 16'hBD15, 16'hD5D8, 16'hDE59, 16'hE69A, 16'hE69B, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE69A, 16'hD619, 16'hDE5A, 16'hE69A, 16'hE65A, 16'hDE59, 16'hDE19, 16'hD597, 16'hC515, 16'hAC52, 16'h9B4E, 16'h930D, 16'hA38F, 16'hBCD4, 16'hD618, 16'hEEDB, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hEEDB, 16'hDDD8, 16'hD598, 16'hE69B, 16'hE65A, 16'hF71D, 16'hFFDF, 16'hDE19, 16'hBC52, 16'hFF5E, 16'hF75E, 16'hDDD9, 16'hF71D, 16'hFFDF, 16'hF71D, 16'hDD98, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hDDD8, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hF71D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF71D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5E,
        16'hFF5E, 16'hFFDF, 16'hFF9F, 16'hCD97, 16'h9C10, 16'hCE18, 16'hDEDB, 16'hD6DA, 16'hD69A, 16'hD69A, 16'hCE18, 16'h4945, 16'hC597, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF
    };

    reg [15:0] image_failed [0:65535] = {
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hEF5D, 16'hDEDB, 16'hD65A, 16'hC618, 16'hBDD7, 16'hB596, 16'h9D13, 16'h9492, 16'h8C51, 16'h8C91, 16'h8C51, 16'h8C51, 16'h9CD3, 16'hA513, 16'hA514, 16'hAD95, 16'hBDD7, 16'hC618, 16'hD69A, 16'hDEDB, 16'hEF9E, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hE71C, 16'hBDD7, 16'hAD55, 16'h9492, 16'h630C, 16'h4208, 16'h3144, 16'h000, 16'h000, 16'h000, 16'h000, 16'h38C2, 16'h730C, 16'h8B8E, 16'h9C50, 16'hA451, 16'hA491, 16'hA451, 16'h9C51, 16'h9410, 16'h8BCF, 16'h8BCF, 16'h838E, 16'h734C, 16'h62CB, 16'h5A8A, 16'h5ACB, 16'h5ACB, 16'h7BCF, 16'h9CD3, 16'hBDD7, 16'hD69A, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hC658, 16'hA514, 16'h7BCF, 16'h5ACA, 16'h3986, 16'h3986, 16'h628A, 16'h730C, 16'h734C, 16'h49C7, 16'h3944, 16'h5A48, 16'h5207, 16'h628A, 16'hB4D3, 16'hD5D7, 16'hDE18, 16'hDE18, 16'hDE18, 16'hDE18, 16'hDE18, 16'hD618, 16'hD618, 16'hD618, 16'hDE18, 16'hDE18, 16'hD618, 16'hD618, 16'hD618, 16'hCDD7,
        16'hC596, 16'hBD55, 16'hACD3, 16'h9410, 16'h7B4D, 16'h62CB, 16'h5A8A, 16'h738E, 16'h8C50, 16'hAD95, 16'hD69A, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hBDD7, 16'h9492, 16'h5ACB, 16'h4A08, 16'h5A8A, 16'h8BCF, 16'hAC92, 16'hBD55, 16'hCD96, 16'hD5D7, 16'hD618, 16'hD618, 16'hD617, 16'hCD96, 16'h838E, 16'h4144, 16'h5A48, 16'hC555, 16'hD618, 16'hD5D7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hCDD7, 16'hB555, 16'hA4D2, 16'h83CF, 16'h62CB, 16'h5ACA, 16'h738E, 16'hA514, 16'hDEDB, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hAD56, 16'h738E, 16'h4A49, 16'h6B0C, 16'h9410, 16'hB514, 16'hCD96, 16'hD618, 16'hD618, 16'hD618, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hCD96, 16'h6A8A, 16'hACD3, 16'hD618, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7,
        16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD618, 16'hD618, 16'hD618, 16'hD658, 16'hD618, 16'hCDD7, 16'hAD14, 16'h8C0F, 16'h5ACB, 16'h4A08, 16'h9492, 16'hCE59, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hEF5D, 16'hE71C, 16'hD69A, 16'hD659, 16'hBD97, 16'hBDD7, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hAD96, 16'h6B4D, 16'h5249, 16'h7B4D, 16'hACD3, 16'hCD96, 16'hD618, 16'hD618, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hD5D7, 16'hC555, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D8, 16'hD618, 16'hD618, 16'hD618, 16'hCE18, 16'hC596, 16'h9C51, 16'h734D, 16'h528A, 16'h9492, 16'hD69A, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hEF5D, 16'hE71C, 16'hD699, 16'hC618, 16'hAD55, 16'h9CD3, 16'h8C10, 16'h738E, 16'h5289, 16'h628B, 16'h628A, 16'h730D, 16'h7B4D, 16'h9C11, 16'h9C11, 16'h83CF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDE, 16'hCE59, 16'h7BCF, 16'h39C7, 16'h734D, 16'hACD3, 16'hCDD7, 16'hD618, 16'hD5D7, 16'hCDD7, 16'hCD97, 16'hCD96, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7,
        16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCD97, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D8, 16'hD5D8, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D8, 16'hD5D8, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D8, 16'hD618, 16'hD618, 16'hD618, 16'hC5D7, 16'h9C92, 16'h6B0C, 16'h5249, 16'h9492, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hE71C, 16'hDEDB, 16'hCE59, 16'hC617, 16'hAD55, 16'h9492, 16'h8C10, 16'h5ACB, 16'h62CB, 16'h5249, 16'h6B0C, 16'h730C, 16'h7B4E, 16'h9C51, 16'hAC93, 16'hC556, 16'hCDD8, 16'hD619, 16'hE65A, 16'hEE9B,
        16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF69C, 16'h838E, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hBDD7, 16'h5ACB, 16'h49C7, 16'h9C51, 16'hC596, 16'hD618, 16'hD5D7, 16'hCDD7, 16'hCD97, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCD97, 16'hCD96, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D8, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D8, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD5D8, 16'hCE17, 16'hCE17, 16'hD618, 16'hD618,
        16'hD618, 16'hBD96, 16'h9450, 16'h4A08, 16'h6B4D, 16'hAD55, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hEF5D, 16'hE71C, 16'hD69A, 16'hC618, 16'hBD96, 16'hAD54, 16'h9CD3, 16'h8C51, 16'h7BCF, 16'h738D, 16'h6B0C, 16'h62CB, 16'h62CB, 16'h7BCF, 16'h8C10, 16'h9C93, 16'hAD14, 16'hBD96, 16'hCDD8, 16'hD659, 16'hE69B, 16'hEEDC, 16'hF71C, 16'hF71C, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hEE9B, 16'hF6DC, 16'hE65A, 16'hCD97, 16'hE619, 16'h7B4D, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hBDD6, 16'h4A49, 16'h6ACB, 16'hB514, 16'hD5D7, 16'hD618, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7,
        16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hC555, 16'hB4D3, 16'hACD3, 16'hACD3, 16'hC555, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD5D8, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hCE18, 16'hCE17, 16'hCE17, 16'hD618, 16'hD659, 16'hCE17, 16'hAD14, 16'h62CB, 16'h630C, 16'hB596, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hEF5D, 16'hDEDB, 16'hCE59, 16'hC618, 16'hAD55, 16'hA4D3, 16'h9492, 16'h8410, 16'h738E, 16'h6B0C, 16'h5ACA, 16'h738D, 16'h734D, 16'h8410, 16'h9C92, 16'hA514, 16'hB556, 16'hC5D7, 16'hD659, 16'hDE9A, 16'hE71C, 16'hF75D, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hF75D, 16'hF71D, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hF6DC, 16'hDE19, 16'h7B0C, 16'hA410, 16'hDD97, 16'h6A8A, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h4A49, 16'h628A, 16'hB514, 16'hD618, 16'hD618, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCD96, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCD97, 16'hC555, 16'hCD96, 16'hC555, 16'hA492, 16'hB4D3, 16'hCD96, 16'hD618, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8,
        16'hD5D8, 16'hD5D8, 16'hD618, 16'hD5D8, 16'hD5D8, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hCE18, 16'hCE17, 16'hCE17, 16'hD618, 16'hD658, 16'hD658, 16'hBD96, 16'h7B8E, 16'h000, 16'h738E, 16'h7B8E, 16'h7BCE, 16'h6B4D, 16'h5289, 16'h5249, 16'h62CB, 16'h83CF, 16'h9451, 16'hA4D3, 16'hB556, 16'hC5D7, 16'hD65A, 16'hE6DB, 16'hF75D, 16'hF75E, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF5D, 16'hF71D, 16'hF71C, 16'hEEDC, 16'hEEDC, 16'hFF1D, 16'hC597, 16'h5A08, 16'hB492, 16'hD555, 16'hD515, 16'h72CB, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h5ACB, 16'h5249,
        16'hB514, 16'hD618, 16'hD618, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCD96, 16'hC555, 16'hC555, 16'hC555, 16'hCD96, 16'hCD97, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D8, 16'hD5D7, 16'hD5D7, 16'hC556, 16'hAC92, 16'h93CF, 16'h9C51, 16'hC555, 16'hD618, 16'hD5D7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hCE18, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hCDD7, 16'hAD14, 16'hACD4, 16'hAD14, 16'hBD96, 16'hD659, 16'hE6DB, 16'hF75D, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hB514, 16'h5187, 16'hBC92, 16'hD515, 16'hCCD4, 16'hCD14, 16'h72CB, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h6B4D, 16'h3945, 16'hACD3, 16'hD618, 16'hD618, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCD96, 16'hBD14, 16'hB4D3, 16'hBD14, 16'hC556, 16'hCD96, 16'hCD97, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D8, 16'hCD97,
        16'hB4D3, 16'h8B8F, 16'h9C11, 16'hCD96, 16'hDE18, 16'hD5D7, 16'hCDD7, 16'hD5D7, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD618, 16'hD618, 16'hD5D8, 16'hD5D8, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hCE18, 16'hD659, 16'hE6DC, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5D, 16'hA493, 16'h61C7, 16'hC493, 16'hD514, 16'hCCD4, 16'hD514, 16'hCCD4, 16'h72CB, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hF79E, 16'hF79E, 16'hF79E, 16'hFF9E, 16'hFF9F, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hF79E, 16'hF79D, 16'hEF5D, 16'hE71C, 16'hDEDB, 16'hD69A,
        16'hCE59, 16'hC618, 16'hC618, 16'hBDD7, 16'hC5D7, 16'hBDD7, 16'h8410, 16'h1840, 16'h9C51, 16'hD617, 16'hD618, 16'hD5D7, 16'hCDD7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hBD55, 16'hAC92, 16'hAC92, 16'hBD55, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD597, 16'hD597, 16'hD5D7, 16'hCDD7, 16'hCD97, 16'hD5D7, 16'hD5D8, 16'hD5D7, 16'hB4D3, 16'h8B8E, 16'hAC92, 16'hD5D8, 16'hD5D8, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hCE18, 16'hDE9A, 16'hEF1D, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'h9410, 16'h6208, 16'hCD14, 16'hD514, 16'hCCD4, 16'hCCD4, 16'hD514, 16'hC493, 16'h730C, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD96, 16'h7B4D, 16'h834D, 16'h730C, 16'h730C, 16'h6ACB, 16'h7B4D, 16'h838E, 16'h7B8D, 16'h7B4E, 16'h7B8E, 16'h7B8E, 16'h83CF, 16'h7BCF, 16'h8410, 16'h840F, 16'h8C10, 16'h8C51, 16'h8C51, 16'h9451, 16'h9492, 16'h9451, 16'h8C51, 16'h9492, 16'h9492, 16'h9451, 16'h9491, 16'h8C51, 16'h9CD2, 16'h8C51, 16'h8C51, 16'h8C51, 16'h7B8E, 16'h840F, 16'h8C10, 16'h738E, 16'h7BCE, 16'h83CF, 16'h738D, 16'h6B4C, 16'h7BCE, 16'h6B4D, 16'h528A, 16'h6B4C, 16'h5ACA, 16'h5289, 16'h5ACA, 16'h5249, 16'h4A08, 16'h4207, 16'h41C7, 16'h5208, 16'h6ACB, 16'h7B4D, 16'h734C, 16'h734D, 16'h4186, 16'h000, 16'h7B4D, 16'hC5D6, 16'hDE58, 16'hD618, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hBD14, 16'hA451, 16'hB4D3, 16'hC596, 16'hD5D7, 16'hD5D8, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7,
        16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD597, 16'hD597, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hD5D8, 16'hCDD7, 16'hA492, 16'h8BCF, 16'hC556, 16'hDE18, 16'hD5D7, 16'hD5D7, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hCE18, 16'hD618, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9E, 16'h7B8E, 16'h728A, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hD514, 16'hBC52, 16'h734D, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h4144, 16'hDDD8, 16'hEE9B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hDE19, 16'hDE59, 16'hD618, 16'hD5D8, 16'hD618, 16'hCD97, 16'hCD97, 16'hC597, 16'hC596, 16'hBD56, 16'hBD96, 16'hB555, 16'hBD55, 16'hBD56, 16'hBD56, 16'hBD56, 16'hBD96, 16'hBD96, 16'hBD96, 16'hBD96, 16'hBDD6, 16'hBDD7, 16'hC5D7, 16'hCE18, 16'hCE18, 16'hCE19, 16'hCE59, 16'hCE18, 16'hCE18, 16'hC5D8, 16'hC5D8,
        16'hBDD7, 16'hC5D7, 16'hC5D7, 16'hBD96, 16'hBD96, 16'hBD55, 16'hBD96, 16'hC5D6, 16'hCDD7, 16'hCE18, 16'hD618, 16'hD618, 16'hDE59, 16'hDE59, 16'hDE99, 16'h9451, 16'h7B8E, 16'hCDD7, 16'hD658, 16'hD618, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hC596, 16'hB4D3, 16'hB4D4, 16'hCD96, 16'hD5D8, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD597, 16'hD597, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hD5D7, 16'hDE18, 16'hC555, 16'h8BCF, 16'hB4D3, 16'hDE18, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hCE18, 16'hD659, 16'hF79E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'h738E, 16'h830C, 16'hD514, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hD515, 16'hB411, 16'h83CF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h4145, 16'hEE9B, 16'hF69C, 16'hF69B, 16'hFF1D, 16'hF6DC, 16'hF6DC, 16'hF71C, 16'hF6DC, 16'hF71C, 16'hF71C, 16'hF71D, 16'hF71D, 16'hFF5D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hEF1C, 16'hE69A, 16'hDE59, 16'hD659, 16'hD618, 16'hD658, 16'hD658, 16'hCE18, 16'hCE18, 16'hCE17, 16'hBD96, 16'hCE18, 16'hD618, 16'hD618, 16'hD5D8, 16'hD5D8, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hCDD7, 16'hCDD7, 16'hD5D8, 16'hD5D7, 16'hC596, 16'hC555, 16'hCDD7, 16'hD618, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hD5D7, 16'hD5D7,
        16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD597, 16'hD597, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCD97, 16'hCD97, 16'hD5D7, 16'hCDD7, 16'h93CF, 16'h9C10, 16'hD618, 16'hD618, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hCE18, 16'hCE18, 16'hEF1C, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'h62CB, 16'h8B0D, 16'hD515,
        16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hDD15, 16'hA38E, 16'h9492, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1D, 16'h4186, 16'hDDD8, 16'hCD56, 16'h7ACC, 16'hCD97, 16'hF71C, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF71C, 16'hF71C, 16'hF71D, 16'hF71D, 16'hFF5D, 16'hF75E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hF75D, 16'hEF1C, 16'hDE9A, 16'hD618, 16'hCE17, 16'hCE18, 16'hCE18, 16'hCE18, 16'hD658, 16'hCE18, 16'hCE18, 16'hD618, 16'hD5D8, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD618, 16'hC596, 16'hC556, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCD97, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCD97, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hD597, 16'hD5D7, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hDE18, 16'hACD3, 16'h8B8E, 16'hD5D7, 16'hD618, 16'hD5D7, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618, 16'hD618,
        16'hCE18, 16'hCE18, 16'hCE18, 16'hD659, 16'hF71C, 16'hFF5D, 16'hF75D, 16'hFF5E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'h628A, 16'h938E, 16'hD515, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hDD15, 16'h930C, 16'hB595, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h62CB, 16'hBCD3, 16'hD555, 16'hAC51, 16'h6208, 16'h93D0, 16'hEE9B, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF71C, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hF75D, 16'hE6DB, 16'hD658, 16'hCE17, 16'hCE18, 16'hCE18, 16'hCE18, 16'hCE18, 16'hCE18, 16'hD617, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD618, 16'hBD54, 16'hB514, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7,
        16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD597, 16'hCD97, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCD97, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCD97, 16'hD5D7, 16'hD597, 16'hCD97, 16'hCD97, 16'hD597, 16'hD5D7, 16'hD5D7, 16'hD5D8, 16'hD5D8, 16'hDE19, 16'hE65A, 16'hE65A, 16'hE69A, 16'hE69B, 16'hE65A, 16'hE69B, 16'hE69B, 16'hE65A, 16'hEE9B, 16'hD5D7, 16'h8B8E, 16'hC596, 16'hDE19, 16'hD5D7, 16'hD618, 16'hD618, 16'hCE18, 16'hCE17, 16'hCE18, 16'hD618, 16'hD618, 16'hDE59, 16'hE69B, 16'hF71D, 16'hFF5D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1D, 16'h62CB, 16'h938E, 16'hD555, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hD515, 16'h7A8A, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h83CF, 16'hB451, 16'hD556, 16'hD515, 16'hCD15, 16'h830D, 16'h624A, 16'hDE18, 16'hFF1D, 16'hEEDC, 16'hF71D, 16'hFF5D, 16'hFF5E, 16'hFF9E, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hDE9A, 16'hCE18, 16'hC617, 16'hCE17, 16'hCE17, 16'hC5D7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hACD3, 16'hBD14, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCDD7, 16'hCD97, 16'hD5D7, 16'hD5D7, 16'hCD96, 16'hD597, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD97, 16'hCD97, 16'hCD96, 16'hCD96, 16'hCD96, 16'hDE18, 16'hDE18, 16'hD597, 16'hD5D8, 16'hDE19, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hEEDC, 16'hEE9B, 16'hE69B, 16'hE69A,
        16'hE65A, 16'hEE9B, 16'hDE19, 16'h93D0, 16'hBD55, 16'hDE19, 16'hD618, 16'hDE59, 16'hE69A, 16'hE69A, 16'hEEDB, 16'hEEDC, 16'hF6DC, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'h5A8A, 16'h9B8E, 16'hD555, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hD4D4, 16'hD4D4, 16'hD514, 16'h6A49, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA4D3, 16'h9B8F, 16'hD556, 16'hCD14, 16'hCD14, 16'hD555, 16'hA410, 16'h3080, 16'hBD55, 16'hFF1D, 16'hFF5D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hF71C, 16'hE69B, 16'hE69A, 16'hE69A, 16'hD659, 16'hCDD8,
        16'hCDD7, 16'hD618, 16'hD5D7, 16'hA451, 16'hB514, 16'hD5D7, 16'hCD97, 16'hCD97, 16'hCDD7, 16'hD5D7, 16'hD618, 16'hDE19, 16'hDE59, 16'hE65A, 16'hE69A, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hDE18, 16'hCD97, 16'hD5D7, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD97, 16'hD5D7, 16'hCD96, 16'hC556, 16'hDDD8, 16'hE65A, 16'hEEDC, 16'hF6DC, 16'hF69C, 16'hEE9B, 16'hDE19, 16'hCD96, 16'hCD96, 16'hE65A, 16'hEE9B, 16'hEEDC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hEE9B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hEE5B, 16'hE65A, 16'h834E, 16'hCD97, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'h5A8A, 16'hAC10, 16'hD555, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hD4D4, 16'hD4D4, 16'hCCD4, 16'h6249, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h728A, 16'hD555, 16'hCD14,
        16'hCD14, 16'hCCD4, 16'hD555, 16'hB493, 16'h4145, 16'hAC93, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hEEDC, 16'hE69A, 16'hD5D7, 16'h9C10, 16'hBD14, 16'hD5D7, 16'hCD97, 16'hD5D8, 16'hDE59, 16'hEE9B, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hF6DC, 16'hDE19, 16'hDDD8, 16'hDE18, 16'hE659, 16'hE65A, 16'hE65A, 16'hDDD8, 16'hD597, 16'hCD56, 16'hD5D8, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1E, 16'hFF1E, 16'hF6DC, 16'hE619, 16'hDE18, 16'hEE9B, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D,
        16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF6DC, 16'hE65A, 16'hE61A, 16'hE61A, 16'hE65A, 16'hE619, 16'h9C11, 16'hEE9B, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1D, 16'h62CB, 16'hAC10, 16'hD515, 16'hCCD4, 16'hCD14, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hD4D4, 16'hD4D4, 16'hD514, 16'hC492, 16'h730C, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDA, 16'h5146, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCCD4, 16'hD515, 16'hC4D4, 16'h51C7, 16'h93D0, 16'hFF5E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hEEDC, 16'h938E, 16'hBD14, 16'hD618, 16'hDE19, 16'hEEDB, 16'hF71C, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hEE9C, 16'hDDD9, 16'hE65A, 16'hF6DC, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hFF1D, 16'hF71D, 16'hF69B, 16'hBD15, 16'hE65A, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hEE9B, 16'hDE19, 16'hE65A, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hEE9B, 16'hE61A, 16'hDE19, 16'hE65A, 16'hE65A, 16'h8B8F, 16'hE65A, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1D, 16'h628B, 16'hAC10, 16'hD555, 16'hCCD4, 16'hCD14, 16'hCD14, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hD4D4, 16'hCCD4, 16'hD515, 16'hAC10, 16'h8C51, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h5208, 16'hBC93, 16'hD515, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hD514, 16'hD555, 16'h830D, 16'h6B0C, 16'hF75D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF6DC, 16'h938F, 16'hC556, 16'hEE9B, 16'hF6DC, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF6DC, 16'hDDD9, 16'hF69C, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hBCD4, 16'hEE9B, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D,
        16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF6DC, 16'hD5D8, 16'hDE5A, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF6DC, 16'hE65A, 16'hE61A, 16'hEE5B, 16'hDE19, 16'h938F, 16'hEE9B, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1D, 16'h5A49, 16'hAC11, 16'hD515, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCD14, 16'hCCD4, 16'hCD14, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hD4D4, 16'hCCD4, 16'hDD15, 16'h934D, 16'hA514,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h7B8F, 16'h9B8F, 16'hD555, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hD514, 16'hD556, 16'h8B4D, 16'h5A4A, 16'hEEDC, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'h8B8F, 16'hD5D8, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hE65A, 16'hF6DC, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF6DC, 16'hBCD4, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hEEDC, 16'hCD97, 16'hEEDC, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hEE9B, 16'hE65A, 16'hEE9C, 16'hD5D8, 16'h8B8F, 16'hF6DD, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D,
        16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'h6ACB, 16'hAC10, 16'hD555, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hCD14, 16'hCD14, 16'hCCD4, 16'hCD14, 16'hCD14, 16'hCCD4, 16'hCCD4, 16'hCCD4, 16'hD4D4, 16'hCCD4, 16'hDD15, 16'h82CB, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h6A09, 16'hD515, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hD514, 16'hCD14, 16'hCD14, 16'hD556, 16'hA3D0, 16'h4186, 16'hDE9A, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'h9C11, 16'hD5D8, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hEE9C, 16'hF6DC, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D,
        16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF6DC, 16'hBCD4, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hE65A, 16'hD5D8, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hEEDC, 16'hE69B, 16'hF6DC, 16'hCD97, 16'hAC52, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'h6B0C, 16'hA3D0, 16'hD555, 16'hCCD4, 16'hCD14, 16'hCCD4, 16'hCD14, 16'hCD14,
        16'hCD14, 16'hCCD4, 16'hCD14, 16'hCD14, 16'hCCD4, 16'hD4D4, 16'hCCD4, 16'hD4D4, 16'hD4D4, 16'hD515, 16'h6A08, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h4105, 16'hCCD4, 16'hD515, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hD514, 16'hCCD4, 16'hCCD4, 16'hDD55, 16'hB451, 16'h3882, 16'hC618, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hBD14, 16'hCD97, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hEE9B, 16'hC515, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hD597, 16'hEE9B, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hEEDC,
        16'hFF1D, 16'hACD3, 16'hB4D4, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF75E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'h838E, 16'hA3CF, 16'hD555, 16'hCCD4, 16'hCD14, 16'hCD14, 16'hCCD4, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCCD4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hCCD4, 16'hD514, 16'hCC93, 16'h6B0C, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h5ACB, 16'hB451, 16'hD515, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCCD4, 16'hD515, 16'hC493, 16'h2800, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hFF1E, 16'hCD97, 16'hC556, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D,
        16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hE65B, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hEE5B, 16'hCD56, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hE65A, 16'hD5D8, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF6DD, 16'hF71D, 16'hA451, 16'hD5D8, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F,
        16'hFFDF, 16'hFF5E, 16'h734D, 16'hA3CF, 16'hDD56, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCCD4, 16'hCCD4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hCCD4, 16'hD515, 16'hB411, 16'h8C51, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9492, 16'h934D, 16'hD515, 16'hCCD4, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hD514,
        16'hCD14, 16'hCCD4, 16'hD515, 16'hC4D3, 16'h5083, 16'hA4D3, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hE65A, 16'hC556, 16'hFF5D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1E, 16'hE65A, 16'hE65B, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hE65A, 16'hD597, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hD597, 16'hEE9C, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D,
        16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hEEDC, 16'h9BD0, 16'hEEDC, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'h83CF, 16'h9B8E, 16'hD556, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCCD4, 16'hCCD4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hCCD4, 16'hD515, 16'h8B0C, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE19, 16'h6208, 16'hD515, 16'hCD14, 16'hD514, 16'hD514, 16'hD514, 16'hD514, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hD515, 16'hD515, 16'h6A08, 16'h8C10, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hCD97,
        16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hFF1E, 16'hEEDC, 16'hCD97, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hFF5E, 16'hDE19, 16'hDDD8, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1E, 16'hE65A, 16'hDE19, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF5E, 16'hDE19, 16'hB4D3, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'h83CF, 16'h9BCF, 16'hDD56, 16'hCCD5, 16'hCD15, 16'hCD14, 16'hCCD4, 16'hCD14, 16'hCD14, 16'hCD14, 16'hD514, 16'hD514, 16'hD514, 16'hD514, 16'hD514, 16'hD514, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD515, 16'h728A, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h4186, 16'hC4D3, 16'hD515, 16'hCD14, 16'hCD14, 16'hCD14, 16'hD514, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hD514, 16'hCCD4, 16'hD515, 16'hD515, 16'h724A, 16'h738D, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hDE19, 16'hEE9B, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hFF5E, 16'hCD97, 16'hE65A, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hFF5E, 16'hDE19, 16'hDDD9, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D,
        16'hFF1D, 16'hFF1D, 16'hF6DC, 16'hD5D8, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF5E, 16'hC515, 16'hD597, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'h9411, 16'h9BCF, 16'hD596, 16'hD515, 16'hD515, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hCD14, 16'hD514, 16'hD514, 16'hD514, 16'hD514, 16'hD514, 16'hD514, 16'hD4D4, 16'hD4D4, 16'hCCD4, 16'hD514, 16'hC493, 16'h730C, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h7B8F, 16'hA3CF, 16'hD515, 16'hCD14, 16'hD514, 16'hCD14, 16'hCD14, 16'hD514, 16'hD514, 16'hD514, 16'hD514, 16'hD4D4, 16'hCCD4, 16'hCCD4, 16'hD4D4, 16'hD555, 16'h8B4D, 16'h5249, 16'hE6DB, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF71D, 16'hEE9B,
        16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hEE9B, 16'hDE5A, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1E, 16'hEE9B, 16'hC515, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hDDD9, 16'hE65A, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hD5D8, 16'hE65B, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF6DC, 16'hAC52, 16'hF6DC, 16'hFF1E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D,
        16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'h9C92, 16'h940F, 16'hDDD7, 16'hC514, 16'hB451, 16'hCD14, 16'hD555, 16'hCD15, 16'hCCD4, 16'hD514, 16'hD514, 16'hCD14, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD514, 16'hD514, 16'hD514, 16'hD4D4, 16'hCCD4, 16'hD515, 16'hB410, 16'h9492, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h7A8A, 16'hD555, 16'hCD14, 16'hD514, 16'hCD14, 16'hCD14, 16'hCD14, 16'hD514, 16'hD514, 16'hD514, 16'hD4D4, 16'hD4D4, 16'hCD14, 16'hCCD4, 16'hD4D4, 16'hD515, 16'hA3D0, 16'h4145, 16'hD65A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'hDE5A, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hE65A, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF5E, 16'hCD97, 16'hDE19, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1E, 16'hDDD8, 16'hE65A, 16'hFF1D,
        16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1E, 16'hE65A, 16'hCD97, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hDE19, 16'hBCD4, 16'hFF1E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hAD14, 16'h8BCF, 16'hDE58, 16'hD5D8, 16'hEEDB, 16'hC596, 16'h8B0D, 16'hA3CF, 16'hCD14, 16'hDD55, 16'hCD14, 16'hCD14, 16'hD514, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD514, 16'hD514, 16'hD514, 16'hD4D4, 16'hCCD4, 16'hD515,
        16'h8B0C, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h59C7, 16'hCD14, 16'hCD14, 16'hCD14, 16'hD514, 16'hD514, 16'hD514, 16'hD514, 16'hD514, 16'hD514, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hCCD4, 16'hDD55, 16'hBC92, 16'h3000, 16'hB595, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD619, 16'hF71C, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hEE9B, 16'hEEDC, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF6DC, 16'hBCD4, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1E, 16'hDDD8, 16'hEE9B, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF6DD, 16'hC515, 16'hF6DD, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1E, 16'hBCD4, 16'hE65A,
        16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hACD3, 16'h8BCF, 16'hDE59, 16'hD659, 16'hEF1C, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hB556, 16'h728A, 16'hABCF, 16'hD515, 16'hD515, 16'hCCD4, 16'hCD14, 16'hD514, 16'hD514, 16'hD514, 16'hD4D4, 16'hD4D4, 16'hD514, 16'hCD14, 16'hD4D4, 16'hD515, 16'h6A8A, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h62CB, 16'hB451, 16'hD515, 16'hCD14, 16'hD514, 16'hD514, 16'hD514, 16'hD514, 16'hD514, 16'hCD14, 16'hD4D4, 16'hCCD4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD515, 16'hCCD4, 16'h724A, 16'h9C92, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE19, 16'hEE9B, 16'hFF1D, 16'hF71D, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hEE9B, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hDDD8, 16'hCD97, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D,
        16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1E, 16'hDDD8, 16'hF69C, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1E, 16'hCD15, 16'hE65A, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF5E, 16'hEE9B, 16'hB4D3, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFEDD, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9E, 16'h9C92, 16'h9C91, 16'hDE59, 16'hDE59, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hE6DC, 16'h9C52, 16'h7A8A,
        16'hBC52, 16'hDD55, 16'hD515, 16'hCD14, 16'hD514, 16'hD514, 16'hD4D4, 16'hD515, 16'hD515, 16'hCD14, 16'hD515, 16'hC452, 16'h7B8E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h7A8B, 16'hD555, 16'hCCD4, 16'hCD14, 16'hCD14, 16'hCCD4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4,
        16'hD4D4, 16'hD4D4, 16'hDD15, 16'hDD55, 16'h7249, 16'h9C92, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE6DB, 16'hDE19, 16'hFF1D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hBD14, 16'hEE9B, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hDE19, 16'hF6DC, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hDDD8, 16'hCD56, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D,
        16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hC515, 16'hDE19, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF75E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h9410, 16'hBD54, 16'hDE99, 16'hD618, 16'hDE59, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h7B0D, 16'h82CB, 16'hC4D3, 16'hD515, 16'hCD14, 16'hD515, 16'hD514, 16'hD514, 16'hD514, 16'hCD14, 16'hD515, 16'h9B4E, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h51C7, 16'hCCD4, 16'hD514, 16'hCD14, 16'hCD14, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hDD55, 16'hBC51, 16'h9C10, 16'hDE18, 16'h9C51, 16'hF75D, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'hCD97, 16'hF71D, 16'hFF1D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hEE9C, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D,
        16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1E, 16'hEE5B, 16'hBD14, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hDE19, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hEE9B, 16'hB492, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF5F, 16'hFF9F, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hFF1E, 16'hEE9B, 16'hBCD4, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1E, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hFF1E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hC5D7, 16'h7B4D, 16'hBD55,
        16'hDE59, 16'hD658, 16'hE69B, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9E, 16'hCDD7, 16'h8B8F, 16'hB452, 16'hD515, 16'hCD14, 16'hD514, 16'hD514, 16'hCD14, 16'hD514, 16'hD515, 16'h6A0A, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h6B4C, 16'hA3D0, 16'hD515,
        16'hCCD4, 16'hD514, 16'hD514, 16'hD514, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hD4D4, 16'hDD15, 16'hABD0, 16'h6ACA, 16'hE6DC, 16'hFFDF, 16'hD618, 16'h8BCF, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hC596, 16'hE65A, 16'hFF1D, 16'hFF1D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1E, 16'hCD56, 16'hDE18, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hDE19, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hBC93, 16'hE65A, 16'hFF5E,
        16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF1D, 16'hF71D, 16'hFF1E, 16'hBCD4, 16'hE65B, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF1D, 16'hF71D, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF6DD, 16'hF71D, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hE69A, 16'h9C51, 16'h9C51, 16'hF71C, 16'hF75E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hE6DB, 16'hEEDB, 16'hEEDB, 16'hEEDB, 16'hF71C, 16'hFF5D, 16'hB514, 16'h934D, 16'hD556, 16'hD515, 16'hD515, 16'hD515, 16'hCD14, 16'hD515, 16'hBC92, 16'h738D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD6, 16'h6A09, 16'hD515, 16'hCCD4, 16'hCD14, 16'hD514, 16'hD514, 16'hD4D4, 16'hD4D4, 16'hD514, 16'hD4D4, 16'hD514, 16'hD4D4, 16'hD4D4, 16'hDD15, 16'h9B4E, 16'h730C, 16'hF71C, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'hA493, 16'hAD14, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE5A, 16'hBD56, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF1D, 16'hEE9B, 16'hF71D,
        16'hF71D, 16'hFF5E, 16'hFF9F, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hB492, 16'hF6DC, 16'hFF1E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hE65A, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hD597, 16'hCD56, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF1D, 16'hF71D, 16'hFF5E, 16'hDE19, 16'hC555, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D,
        16'hF71D, 16'hFF1D, 16'hEE9C, 16'hF71D, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hF71D, 16'hEEDB, 16'hE69A, 16'hEE9B, 16'hEEDB, 16'h9410, 16'hAD13, 16'hDE9A, 16'hE69A, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hEF1C, 16'hD618, 16'hD5D7, 16'hDE18, 16'hBD55, 16'h7B4D, 16'h834D, 16'hCD15, 16'hD515, 16'hD515, 16'hD515, 16'hCD15, 16'hCD14, 16'hD556, 16'h9B8E, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h4187, 16'hBC93, 16'hD515, 16'hCD14, 16'hD514, 16'hD514, 16'hD514, 16'hD514, 16'hD514, 16'hD4D4, 16'hD514, 16'hCCD4, 16'hDD15, 16'h934E, 16'h7B8E, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hBD56, 16'h8BCF, 16'hE6DB, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'hA452, 16'hF6DC, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1E, 16'hFF1E, 16'hFF1D, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1E, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1E, 16'hE61A, 16'hB4D3, 16'hFF1E, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hE65A, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D,
        16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hEE5A, 16'hBC93, 16'hFF1E, 16'hF71D, 16'hFF5E, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hBCD4, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hE65A, 16'hE69B, 16'hD618, 16'hDE59, 16'hE65A, 16'hDE59, 16'hD5D7, 16'hBD14, 16'h9410, 16'h8BCE, 16'hBD96, 16'hDE9A, 16'hE6DB, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hCE18, 16'hA452, 16'hA492, 16'hB492, 16'hD556, 16'hD555, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hCD15, 16'hD515, 16'h6A49, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9CD2, 16'h8B0C, 16'hD555, 16'hCD14, 16'hD514, 16'hD514, 16'hD515, 16'hD514, 16'hD514, 16'hD514, 16'hD4D4, 16'hDD15, 16'hABD0, 16'h6B0C, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9E, 16'hE69A, 16'hE69A, 16'hD659, 16'h9410, 16'hCDD8, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hB514, 16'hD5D8, 16'hFF5E, 16'hF71D,
        16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF6DC, 16'hF6DD, 16'hF71D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hF71D, 16'hFF5E, 16'hFF9F, 16'hFF1E, 16'hF71D, 16'hFF5E, 16'hF71D, 16'hF6DD, 16'hF71D, 16'hFF5E, 16'hC555, 16'hCD97, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF6DD, 16'hEE9B, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hFEDD, 16'hBC92, 16'hF6DC, 16'hFF1E, 16'hFF5F, 16'hFF9F, 16'hFF5E, 16'hF71D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF5E, 16'hD5D7, 16'hD5D8, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D,
        16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hEE9C, 16'hCD56, 16'hB4D3, 16'h9C51, 16'h9C51, 16'h8BCE, 16'h8BCF, 16'hA451, 16'hCD96, 16'hEEDC, 16'hFF5E, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hAD14, 16'hA410, 16'hDDD7, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hCD15, 16'hD555, 16'hBC52, 16'h734D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71B, 16'h4986, 16'hCD15, 16'hD515, 16'hCD14, 16'hD515, 16'hD515, 16'hCD14, 16'hD515, 16'hD514, 16'hDD15, 16'hB451, 16'h628A, 16'hF71D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hD659, 16'hD618, 16'hC596, 16'hCE17, 16'h7B0C, 16'hBD56, 16'hFF5E, 16'hFFDF, 16'hDE5A, 16'h9410, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hEE9B, 16'hE69B, 16'hFF1D, 16'hF71D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hF71D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF1E, 16'hFF5E, 16'hFF9F, 16'hFF5E, 16'hF6DD, 16'hF71D, 16'hFF1E, 16'hAC92, 16'hEE5B, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hFF1E, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E,
        16'hF6DD, 16'hEE9B, 16'hFF1E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF1E, 16'hC4D4, 16'hE65A, 16'hFF5E, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hEEDC, 16'hC556, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hDDD9, 16'hD618, 16'hDE58, 16'hC5D6, 16'hCDD7, 16'hD618, 16'hEEDB, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hAD14, 16'h6A49, 16'hD556, 16'hD555, 16'hD555, 16'hD555, 16'hD515, 16'hCD14,
        16'hD556, 16'h8B0D, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h83CF, 16'h9BD0, 16'hD555, 16'hCD14, 16'hD515, 16'hD515, 16'hCD15, 16'hD515, 16'hD515, 16'hCD14, 16'h8B4D, 16'hE6DC, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hDE5A,
        16'hDE59, 16'h838E, 16'h734C, 16'hCD97, 16'hBD15, 16'hEF1D, 16'hFF9F, 16'h8BCF, 16'hDE19, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1E, 16'hCD56, 16'hE69B, 16'hFF1D, 16'hF71D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hFF1E, 16'hFF9F, 16'hFF5E, 16'hF71D, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hF6DD, 16'hFF1E, 16'hEE9B, 16'hA451, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hFF9F, 16'hFF5F, 16'hFF1E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hF6DD, 16'hF6DC, 16'hFF1E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF1E, 16'hD597, 16'hD597, 16'hFF5E, 16'hFF1E, 16'hFF5F, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D,
        16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hCD97, 16'hEE9B, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF6DC, 16'hC515, 16'hD618, 16'hD618, 16'hCDD7, 16'hDE59, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hB515, 16'h830D, 16'hD556, 16'hD555, 16'hD555, 16'hD515, 16'hD515, 16'hCD15, 16'h6249, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h51C6, 16'hD555, 16'hD515, 16'hD515, 16'hD515, 16'hD515, 16'hCD15, 16'hD555, 16'hABD0, 16'hAC92, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF75D, 16'hDE59, 16'hDE59, 16'h9C92, 16'hACD3, 16'hE69A, 16'hFF9F, 16'hBD56, 16'h9C51, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hEE9B, 16'hB4D4, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF5E, 16'hFF9F, 16'hFF5E, 16'hF71D, 16'hFF5E, 16'hD5D8, 16'hBD15, 16'hFF5E, 16'hF6DD, 16'hFF1D, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF6DC, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF1E, 16'hE65A, 16'hBCD4, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hE65A, 16'hE65A, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1E, 16'hCD56, 16'hCDD7, 16'hE6DB, 16'hE69B, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hA493, 16'h9B8E, 16'hDD96, 16'hD555, 16'hCD15, 16'hD556, 16'hA410, 16'h8410, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h6B4C, 16'hAC51, 16'hD556, 16'hCD15, 16'hCD15, 16'hCD15, 16'hCD15, 16'hD555,
        16'hCD15, 16'h9BCF, 16'h6A8B, 16'hBD56, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF71D, 16'hDE5A, 16'hDE59, 16'h9C51, 16'hAC92, 16'hDE59, 16'h730C, 16'hE69B, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF6DD, 16'hFF1E, 16'hC556, 16'hD598, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF5E, 16'hBCD4, 16'hD5D8, 16'hFF5E, 16'hF6DD, 16'hF71D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF6DD, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF9F, 16'hFF5E, 16'hFF1D, 16'hF6DC, 16'hB452, 16'hF6DD, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D,
        16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF6DD, 16'hDE19, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hE65A, 16'hB4D3, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1D, 16'hA4D4, 16'h7B4D, 16'hBCD3, 16'hD555, 16'hD555, 16'hD515, 16'hD556, 16'h6209, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h6A49, 16'hD556, 16'hCD15, 16'hCD15, 16'hD515, 16'hD555, 16'hD555, 16'hD555, 16'hDD96, 16'hCD14, 16'h82CB, 16'h730C, 16'hD65A, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hEEDB, 16'hBD55, 16'hD5D7, 16'h9C51, 16'hA452, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF6DC, 16'hAC52, 16'hF6DC, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D,
        16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hAC51, 16'hEE9B, 16'hFF1E, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF9F, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF6DD, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hC4D4, 16'hE65A, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hDE19, 16'hF6DC, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hB493, 16'hCDD8,
        16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF75E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF75E, 16'hDE9A, 16'hA493, 16'h7B0C, 16'h93CF, 16'hCD55, 16'hD556, 16'hD555, 16'hD555, 16'hD556, 16'hC4D3, 16'h62CA, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h5A89, 16'hB493, 16'hD556, 16'hD515, 16'hD515, 16'hD555, 16'hD555, 16'hD555, 16'hD555, 16'hD556, 16'hDD97, 16'hC514, 16'h8B4D, 16'hBD55, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hE6DB, 16'hD618, 16'hCDD7, 16'h6289, 16'hE69B, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1E, 16'hD5D8, 16'hBD15, 16'hFF1E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF6DC, 16'hA411, 16'hF6DD, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D,
        16'hFF1D, 16'hF71D, 16'hFF5E, 16'hD556, 16'hD597, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1E, 16'hDE19, 16'hE65A, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1E, 16'hDDD9, 16'h8B8D, 16'hD618, 16'hE69A, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hEEDC, 16'hC556, 16'hF6DC, 16'hE65A, 16'hE659, 16'hB4D4, 16'h9BCF, 16'hAC51, 16'hCD55, 16'hD596, 16'hD556, 16'hD555, 16'hD556, 16'hD555, 16'hDD96, 16'h8B4D, 16'hA554, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD96, 16'h6209, 16'hD556, 16'hD555, 16'hD555, 16'hD555, 16'hD555, 16'hD555, 16'hD556, 16'hD556, 16'hD556, 16'hDD97, 16'hD597, 16'hCD55, 16'hE69B, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hEEDC, 16'hCDD7, 16'hDE59, 16'h9C10, 16'hAC93, 16'hFF5E, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hAC93, 16'hE65A,
        16'hFF1E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hEE5B, 16'hAC52, 16'hFF1E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hE619, 16'hC4D4, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hEE9B, 16'hD5D8, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D,
        16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'h93CF, 16'hC555, 16'hCDD7, 16'hD618, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hBD96, 16'hAC51, 16'hDD97, 16'hCD55, 16'hD556, 16'hDD97, 16'hDD96, 16'hD556, 16'hCD55, 16'hCD55, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'h5A08, 16'hDF1C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h5ACA, 16'hB493, 16'hD596, 16'hD555, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD596, 16'hCD56, 16'hDE18, 16'hD5D8, 16'hE69B, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF71C, 16'hCDD7, 16'h5A08, 16'hE69B, 16'hFF1D, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1E, 16'hEE5B, 16'hA451, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hDDD8, 16'hB493, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D,
        16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hEE9C, 16'hBC93, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF6DC, 16'hC556, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hFF1D, 16'hBD15, 16'h9C51, 16'hEE9B, 16'hE6DB, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'h8BD0, 16'hC514, 16'hD596, 16'hCD55, 16'hCD55, 16'hCD55, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD555, 16'hDD96, 16'hAC52, 16'h7BCF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC5D8, 16'h5207, 16'hD596, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hDDD8, 16'hBD14, 16'h9BD0, 16'hF71D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hEEDB, 16'h9C10, 16'h9C51, 16'hFF5E, 16'hF71D, 16'hFF1D,
        16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF5E, 16'hBD15, 16'hCD96, 16'hFF5E, 16'hF6DD, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hCD56, 16'hC556, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hB493, 16'hF6DC, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D,
        16'hC556, 16'hE65A, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hE61A, 16'h834D, 16'hDE59, 16'hF71D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE69B, 16'h830D, 16'hD596, 16'hCD55, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hDD97, 16'h6A8A, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h6B4D, 16'hAC92, 16'hDD97, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hDDD7, 16'hB492, 16'h730C, 16'hEF1C, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hE69B, 16'hD618, 16'h5A08, 16'hDE59, 16'hFF5D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hA411, 16'hEE9B, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hBCD4, 16'hD5D7, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D,
        16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hBC93, 16'hE65A, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hDDD8, 16'hD5D8, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'h9C11, 16'hBD55, 16'hF75D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'h9451, 16'hAC51, 16'hD596, 16'hCD55, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556,
        16'hDD97, 16'hC4D4, 16'h6B0C, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h59C8, 16'hD596, 16'hD556, 16'hD596, 16'hD556, 16'hD556, 16'hD556, 16'hDDD7, 16'hAC51, 16'h6B0C, 16'hF71D, 16'hFFDF,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hE69B, 16'hE65A, 16'hACD3, 16'h8BCF, 16'hFF5D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1E, 16'hE65A, 16'hA451, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hBC93, 16'hDE19, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hC515, 16'hDDD8, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D,
        16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hE65A, 16'hBD15, 16'hFF1E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFEDD, 16'hC556, 16'hACD3, 16'hFF5E, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE69B, 16'h6A8A, 16'hCD96, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hD556, 16'hDD97, 16'h728A, 16'hB5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h7B8E, 16'hA452, 16'hD5D7, 16'hD596, 16'hD596, 16'hD596, 16'hD597, 16'hAC52, 16'h7B4E, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hEEDC, 16'hDE19, 16'hE65A, 16'h730C, 16'hD5D8, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF6DD, 16'hFF5E, 16'hC515, 16'hC556, 16'hFF1E, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hB452, 16'hE65A, 16'hFF5E,
        16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hD5D8, 16'hC515, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF6DD, 16'hEE9B, 16'hBD15, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hFF1D, 16'hFF5E, 16'hE69B, 16'hCDD8, 16'hCDD8, 16'hE69B, 16'hFF1D, 16'hF6DD, 16'hF71D, 16'hE61A, 16'h93CF, 16'hC596, 16'hA451, 16'hB555, 16'hE6DB, 16'hFF9E, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB555, 16'h93CF, 16'hD597, 16'hD556, 16'hD596, 16'hD596, 16'hD596, 16'hDD97, 16'hC514, 16'h630B, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hDEDA, 16'h49C7, 16'hCD96, 16'hD596, 16'hD596, 16'hD596, 16'hD596, 16'h7B0C, 16'h83CF, 16'hCE19, 16'hEF1C, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'hDE59, 16'hE659, 16'hC556, 16'h7B4D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hA410, 16'hE65A, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hAC11, 16'hEE9B, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hE61A, 16'hB452, 16'hFF1E, 16'hF71D,
        16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hEE9B, 16'hB4D4, 16'hEE9B, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF5E, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hFF1E, 16'hEEDC, 16'h9C52, 16'h528A, 16'h634E, 16'h73D0, 16'h5ACB, 16'hD619, 16'hFF1D, 16'hF71D, 16'hF6DC, 16'hAC52, 16'hB513, 16'hD5D7, 16'h9C10, 16'h6ACB, 16'h7B4D, 16'h9451, 16'hAD55, 16'hC5D7, 16'hC5D8, 16'hCE18, 16'hAD14, 16'h6A49, 16'hD596, 16'hD596, 16'hD596, 16'hD596, 16'hD556, 16'hDDD7, 16'h8B8E, 16'h528A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9451, 16'h93CF, 16'hD5D7, 16'hCD96, 16'hD596, 16'hD596, 16'hD597, 16'hBCD4, 16'h834D, 16'h730C, 16'h7B8E, 16'h8C10, 16'hA4D3, 16'h9411, 16'h8BCF, 16'hC555, 16'h8B8E, 16'hBD55, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hEE9B, 16'hA411, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D,
        16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFEDD, 16'hAC11, 16'hF6DC, 16'hFF1E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hF69C, 16'hAC51, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hBD15, 16'hDE19, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hCD97, 16'h9C52, 16'hACD4, 16'hCD97, 16'hF6DC, 16'hFF1E, 16'hFF1D, 16'hDE5A, 16'h62CB, 16'h7C10, 16'hADD7, 16'hADD8, 16'hB619,
        16'h8492, 16'h8BD0, 16'hFF1D, 16'hF6DC, 16'hF6DC, 16'hD5D7, 16'h8BCF, 16'hDE18, 16'hD5D8, 16'hD597, 16'hBD15, 16'hAC92, 16'h93CF, 16'h8B8E, 16'h93CF, 16'h9410, 16'h9C51, 16'hBCD4, 16'hD596, 16'hD596, 16'hD596, 16'hD596, 16'hD596, 16'hC555, 16'h4A08, 16'h3985, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h41C7, 16'hC555, 16'hD5D7, 16'hD597, 16'hD597, 16'hD597, 16'hD5D7, 16'hDDD7, 16'hD597, 16'hC515, 16'hBD14, 16'hB4D3, 16'hBD14, 16'hCD97, 16'hC555, 16'h6A8A, 16'hEEDB, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF6DD, 16'hFF5E, 16'hCD97, 16'hBD15, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF6DC, 16'hA3D0, 16'hF6DC, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D,
        16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hF6DD, 16'hA410, 16'hF6DC, 16'hFF1E, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hC515, 16'hCD97, 16'hFF5E, 16'hF6DD, 16'hFF1E, 16'hB515, 16'h3A89, 16'h8CD3, 16'h8493, 16'h5B4D, 16'h5ACB, 16'hC597, 16'hEEDC, 16'h524A, 16'h8CD3, 16'hBE19, 16'hADD8, 16'hADD8, 16'hADD8, 16'h9D15, 16'h734E, 16'hF6DC, 16'hF6DD, 16'hF6DC, 16'hE61A, 16'h8B8F, 16'hC595, 16'hD597, 16'hCD97, 16'hD5D7, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hD5D8, 16'hC556, 16'hC555, 16'hDE18, 16'hD5D7, 16'hD596, 16'hD596, 16'hCD96, 16'hD5D7, 16'h8B8E, 16'h7B4E, 16'hACD3, 16'h6B4C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB595, 16'h730C, 16'hD5D7, 16'hD597, 16'hD597, 16'hD597, 16'hD597, 16'hD596, 16'hD597, 16'hD5D7, 16'hD5D7, 16'hDE18, 16'hD5D7, 16'hDE18, 16'h8B8E, 16'hA492, 16'hFF1D, 16'hF71C, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF1E, 16'hB4D3,
        16'hD5D8, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF69C, 16'hABD0, 16'hF6DC, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hAC11, 16'hE65A, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hEE9B, 16'hF6DC, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hFF1D, 16'hCD57, 16'hB4D4, 16'hFF5E, 16'hFF1D, 16'hF6DC, 16'h630C, 16'hA5D7,
        16'hB619, 16'hAE19, 16'hAE19, 16'h9555, 16'h5B0C, 16'h41C6, 16'h8452, 16'hB619, 16'hA5D8, 16'hADD8, 16'hADD8, 16'hADD8, 16'hA556, 16'h6B0C, 16'hEEDB, 16'hF71D, 16'hF6DD, 16'hEE9B, 16'h9C10, 16'hA451, 16'hD5D8, 16'hCD97, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hC556, 16'h93D0, 16'h8BCF, 16'hD5D7, 16'hD5D7, 16'hCD96, 16'hD597, 16'hCD55, 16'h4186, 16'hB514, 16'hD5D8, 16'h62CB, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h5249, 16'hACD3, 16'hD5D8, 16'hCD97, 16'hD5D7, 16'hD5D7, 16'hD597, 16'hCD96, 16'hD597, 16'hD5D7, 16'hCD97, 16'hD5D7, 16'hCD96, 16'h5A49, 16'hE65A, 16'hF71D, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hFF1D, 16'hF6DC, 16'hA411, 16'hEE9B, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF69C, 16'hAC11, 16'hF6DD, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D,
        16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF5E, 16'hB492, 16'hDDD9, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hE65B, 16'hEE9B, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hFF1D, 16'hE619, 16'h9C11, 16'hF71D, 16'hFF1E, 16'hDE1A, 16'h5B0C, 16'hADD8, 16'hA598, 16'hA5D7, 16'hA597, 16'hADD8, 16'hA5D7, 16'h7C52, 16'hA5D8, 16'hA5D8, 16'hA5D8, 16'hADD8, 16'hADD8, 16'hADD8, 16'hAD97, 16'h6B4D, 16'hEEDB, 16'hF71D, 16'hF6DD, 16'hF6DC, 16'hBD15, 16'h8B8E, 16'hD5D7, 16'hCD97, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD97, 16'hD5D7, 16'hA451, 16'h7B4D, 16'hD5D7, 16'hD5D6, 16'hD5D7, 16'h8B8F, 16'h6B0D, 16'hCDD7, 16'hD5D7, 16'hACD3, 16'h7BCE, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE58, 16'h4186, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD597, 16'hCD96, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D8, 16'h9410, 16'h838E, 16'hF71D, 16'hF6DD, 16'hF71D,
        16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hFF1E, 16'hE65A, 16'hAC52, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hF69C, 16'hAC11, 16'hF6DD, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF5E, 16'hBCD4, 16'hCD56, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hEE9B, 16'hE65A,
        16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DC, 16'hF71D, 16'hEE9B, 16'h938F, 16'hEE9B, 16'hFF1D, 16'hEE9B, 16'h5ACC, 16'hA5D7, 16'hA5D8, 16'hADD8, 16'hAE19, 16'hAE18, 16'hADD8, 16'hA5D8, 16'hA5D7, 16'hA5D8, 16'hADD8, 16'hADD8, 16'h9515, 16'hA596, 16'h94D4, 16'h838F, 16'hFF1D, 16'hF71C, 16'hF71D, 16'hF6DC, 16'hD597, 16'h7B4D, 16'hCD96, 16'hCD97, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hDE59, 16'hACD3, 16'h7B4D, 16'hD5D7, 16'hBD14, 16'h3145, 16'hBD55, 16'hCDD7, 16'hCD96, 16'hCDD7, 16'h5208, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h8410, 16'h9410, 16'hDE18, 16'hCD97, 16'hCDD7, 16'hCD97, 16'hCD96, 16'hC555, 16'hC555, 16'hC555, 16'hC596, 16'h49C7, 16'hC597, 16'hF71D, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hCD97, 16'hBD14, 16'hF71D, 16'hF6DC, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hEE5B, 16'hB452, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D,
        16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hFF5E, 16'hC556, 16'hB492, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hEE9B, 16'hDE19, 16'hF6DD, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'h93D0, 16'hDE1A, 16'hFF1E, 16'hF6DC, 16'h738E, 16'hA5D7, 16'hB619, 16'hA596, 16'h8493, 16'h8CD4, 16'hA597, 16'hADD8, 16'h9D97, 16'hADD8, 16'h9515, 16'h5ACC, 16'h830D, 16'h834E, 16'h5A49, 16'h630C, 16'hDE9A, 16'hFF1D, 16'hF6DD, 16'hF6DD, 16'hE65A, 16'h93CF, 16'hB4D4, 16'hD5D7, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD97, 16'hCD97, 16'hACD3, 16'h838E, 16'h83CE,
        16'hD596, 16'h628A, 16'h9451, 16'hCDD7, 16'hCD96, 16'hCD97, 16'hD5D8, 16'h9C11, 16'h9492, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h3986, 16'hBD54, 16'hD618,
        16'hACD3, 16'h8BCF, 16'h9C51, 16'h9410, 16'h9C51, 16'hA492, 16'h838E, 16'h62CB, 16'hEEDC, 16'hEEDC, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1E, 16'hB4D4, 16'hCD97, 16'hF71D, 16'hF6DC, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hEE5B, 16'hB452, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF6DD, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF6DD, 16'hFF1E, 16'hD5D8, 16'h9C10, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD,
        16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF71D, 16'hEE9B, 16'hDDD8, 16'hF6DC, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hFF1D, 16'hA492, 16'hC597, 16'hFF1E, 16'hFF1D, 16'h9410, 16'h84D3, 16'h7411, 16'h5A8A, 16'h9C10, 16'hA411, 16'h62CB, 16'h8452, 16'hADD8, 16'h9555, 16'h62CB, 16'hCCD5, 16'hFE19, 16'hF5D8, 16'hE597, 16'hD516, 16'h830D, 16'hB515, 16'hFF1D, 16'hF6DD, 16'hF6DC, 16'hB493, 16'h93D0, 16'hD5D7, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD97, 16'hD597, 16'hBD14, 16'h9410, 16'h9C51, 16'hB514, 16'hC596, 16'h8B8F, 16'h6ACB, 16'hCDD7, 16'hCD97, 16'hCD97, 16'hD5D7, 16'hD5D7, 16'hCD97, 16'h5A8A, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h5249, 16'hD618, 16'hC596, 16'h9410, 16'h9C51, 16'hC596, 16'hC596, 16'hDE18, 16'h6ACB, 16'hB514, 16'hF71D, 16'hEEDC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hAC52, 16'hE65A, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF6DD, 16'hFF1E,
        16'hEE5A, 16'hB452, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hEE9C, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hFF1E, 16'hE65A, 16'h834D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF69C, 16'hDDD8, 16'hEE9B, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hFF1D, 16'hBD15, 16'hB4D5, 16'hFF1D, 16'hFF1D, 16'hCD97, 16'h000, 16'hAC11, 16'hEDD9, 16'hFE1A, 16'hF619, 16'hE597, 16'h7A8B, 16'h7C11, 16'h63CF, 16'hAC11, 16'hFE5A, 16'hF5D8, 16'hF5D9, 16'hFE19, 16'hFE5A, 16'hFE1A, 16'h7ACC, 16'hCDD7, 16'hFF1D, 16'hF6DC, 16'hC556,
        16'h7B0C, 16'hD597, 16'hCD97, 16'hCD96, 16'hCD96, 16'hCD96, 16'hA492, 16'hACD3, 16'hC556, 16'hD5D7, 16'hD5D7, 16'hB4D3, 16'h5209, 16'hBD55, 16'hCDD7, 16'hCD96, 16'hCD97, 16'hCDD7, 16'hCDD7, 16'hDE18, 16'h7B4D, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h6B4C, 16'hA492, 16'hDE18, 16'hD618, 16'hB514, 16'h9C51, 16'hAC92, 16'hB514, 16'h5208, 16'hE69A, 16'hF71C, 16'hF71C, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hEE9C, 16'hA411, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF6DD, 16'hFF1D, 16'hEE5A, 16'hBC52, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hEE9B, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD,
        16'hFF1D, 16'hEE9B, 16'h6A8A, 16'hEE9B, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hDDD8, 16'hE65A, 16'hF71D, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hFF1D, 16'hCD97, 16'h9C52, 16'hFF1D, 16'hF6DC, 16'h7B4D, 16'hBC93, 16'hFE1A, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hFE1A, 16'hED98, 16'h6A4B, 16'h4208, 16'hDD56, 16'hED97, 16'hCC93, 16'hDD15, 16'hFE19, 16'hF5D9, 16'hFE5A, 16'hCD15, 16'h9451, 16'hFF1D, 16'hF6DC, 16'hDE18, 16'h7B0C, 16'hC555, 16'hD5D7, 16'hCD96, 16'hCD96, 16'hCD97, 16'hA492, 16'h838E, 16'hB514, 16'hB514, 16'hB4D3, 16'hC555, 16'h9410, 16'h9410, 16'hCDD7, 16'hCD96, 16'hCD96, 16'hCDD7, 16'hCDD7, 16'hD5D8, 16'hBD55, 16'h62CB, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h4186, 16'hC596, 16'hD618, 16'hDE19, 16'hC596, 16'hBD55, 16'h838E, 16'h9410, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hDE19, 16'hB493, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D,
        16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF6DD, 16'hF6DC, 16'hFF1D, 16'hEE5A, 16'hB411, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hE65B, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF6DD, 16'hFF1D, 16'hEE9B, 16'h59C7, 16'hE65A, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hDDD8, 16'hE659, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hDE19, 16'h8BCF, 16'hFF1D, 16'hACD3, 16'hAC11, 16'hFE1A, 16'hF5D9, 16'hF5D9, 16'hED98, 16'hDD56, 16'hE557, 16'hFE19, 16'hBC93, 16'h1800,
        16'hCCD4, 16'hCC93, 16'hC452, 16'hDD15, 16'hFE19, 16'hF5D9, 16'hFE1A, 16'hD515, 16'h9411, 16'hFF1D, 16'hF6DC, 16'hEE5B, 16'h938F, 16'hB4D3, 16'hD5D7, 16'hCD96, 16'hC555, 16'hACD3, 16'hD5D7, 16'hAC92, 16'h7B4E, 16'hB514, 16'h8C0F, 16'h7B4D, 16'h93D0, 16'hBD14, 16'hCD97, 16'hCD96, 16'hCD96, 16'hCD97, 16'hD5D7, 16'hCDD7, 16'hD5D7, 16'h628A, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h6ACB, 16'hD618, 16'hBD15, 16'hB4D4, 16'hCD96, 16'h5A49, 16'hCDD7, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hFF1E, 16'hCD57, 16'hC515, 16'hF6DD, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hFF1D, 16'hEE5A, 16'hAC11, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D,
        16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hE65B, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hFF1D, 16'hEE9B, 16'h4104, 16'hCD97, 16'hFF1D, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hDDD9, 16'hDE19, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hF6DC, 16'hE65A, 16'h8B8F, 16'hE65B, 16'h834E, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hC493, 16'hABCF, 16'hA38E, 16'hABD0, 16'h9B8F, 16'h628A, 16'hCCD4, 16'hCCD4, 16'hDD16, 16'hF5D8, 16'hF5D9, 16'hF5D9, 16'hFE1A, 16'hAC11, 16'hA4D4, 16'hFF1D, 16'hF6DC, 16'hF6DC, 16'hAC92, 16'h93CF, 16'hD5D7, 16'hCD96, 16'hCD96, 16'hB514, 16'h8BCF, 16'h9410, 16'h730C, 16'hCD96, 16'hD5D7, 16'hCD96, 16'hCD97, 16'hCD97, 16'hCD96, 16'hCD97, 16'hCD96, 16'hCD96, 16'hD5D7, 16'hCDD7, 16'hD5D8, 16'hA492, 16'h8C51, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9451, 16'hACD3, 16'hACD3, 16'hBD55, 16'hB4D3, 16'h628B, 16'hEEDB, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF6DC,
        16'hFF1D, 16'hC4D4, 16'hD597, 16'hF6DD, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hEE5A, 16'hABD1, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hEE5B, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hF6DD, 16'hEE9B, 16'h4083, 16'hB4D4, 16'hFF1D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hDE19, 16'hDDD8, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEEDC, 16'hF69B, 16'h9C11,
        16'hC556, 16'h9B90, 16'hFE19, 16'hF5D9, 16'hF5D9, 16'hF619, 16'hCCD4, 16'hAC11, 16'hC453, 16'hE557, 16'hCCD5, 16'h000, 16'hDD56, 16'hFE19, 16'hF5D9, 16'hF5D8, 16'hF5D8, 16'hF5D9, 16'hF5D9, 16'h6A8A, 16'hD619, 16'hFF1D, 16'hF6DC, 16'hF6DC, 16'hD597, 16'h7B0C, 16'hCD97, 16'hCD96, 16'hCD96, 16'hCDD7, 16'hC596, 16'h9C10, 16'hA492, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD56, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD97, 16'hBD55, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hC596, 16'h5A8A, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h5A48, 16'hB514, 16'hC596, 16'h838D, 16'hA492, 16'hF6DC, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hB452, 16'hDE19, 16'hF6DD, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DD, 16'hEE5A, 16'hA3D0, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D,
        16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hEE5B, 16'hF6DC, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hEE9C, 16'h4946, 16'h9BD0, 16'hFEDD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hE619, 16'hDDD8, 16'hEE9B, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hA452, 16'hBCD5, 16'h9BD0, 16'hF619, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hFDD9, 16'hFE1A, 16'hB452, 16'h0C3, 16'h6A8A, 16'hDD56, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hEDD8, 16'h830D, 16'h9C52, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hDE19, 16'h72CB, 16'hC556, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD97, 16'hCDD7, 16'hCD97, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD97, 16'hC555, 16'hC556, 16'hD5D7,
        16'hCDD7, 16'hD618, 16'h730C, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC5D7, 16'h4185, 16'hB514, 16'h3945, 16'hCDD7, 16'hEEDB, 16'hEE9B,
        16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hEEDC, 16'hBCD3, 16'hEE5B, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hEE9C, 16'hF6DC, 16'hF6DC, 16'hEE1A, 16'h9B8F, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hEE5B, 16'hEE9C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF69C, 16'h6249, 16'h72CB, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC,
        16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hE619, 16'hD597, 16'hEE5B, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DD, 16'hB4D4, 16'hC556, 16'h8BD0, 16'hD515, 16'hFE1A, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hF5D9, 16'hFDD9, 16'hE597, 16'h5209, 16'h7C50, 16'h5B0C, 16'h4A08, 16'h834D, 16'h9BCF, 16'h830C, 16'h5248, 16'h1144, 16'hA493, 16'hFF1D, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hEE9B, 16'h7ACC, 16'hB4D3, 16'hCDD7, 16'hCD96, 16'hCD96, 16'hCD96, 16'hC556, 16'hDE59, 16'hDE59, 16'hC555, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hB514, 16'hD5D7, 16'hD5D7, 16'hD618, 16'hB514, 16'h6B4D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9C93, 16'h000, 16'h734D, 16'hEEDB, 16'hE69A, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hEE5A, 16'hC515, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hEE5A, 16'h9B8F, 16'hEEDC, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF71D,
        16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hEE5B, 16'hEE9C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'h7ACC, 16'h4945, 16'hEE9B, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hDE19, 16'hD597, 16'hEE5A, 16'hEEDC, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hF6DD, 16'hB4D4, 16'hB4D4, 16'hD619, 16'h3903, 16'hD516, 16'hFE1A, 16'hFE1A, 16'hFE19, 16'hFE1A, 16'hEDD8, 16'h728A, 16'h7C50, 16'h9514, 16'h8492, 16'h9D14, 16'h8C51, 16'h8C51, 16'h9492, 16'h94D3, 16'hAD96, 16'h3186, 16'hDE19, 16'hFF1D, 16'hF6DC, 16'hF71C, 16'hF6DC, 16'h9BD0, 16'h9C51, 16'hD5D7, 16'hC596, 16'hCD96, 16'hC556, 16'hCD97,
        16'hEEDC, 16'hF6DC, 16'hCDD7, 16'hC556, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hD5D7, 16'hB514, 16'hCD96, 16'hD5D8, 16'hD5D7, 16'hD5D8, 16'h62CB, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h62CB, 16'hA493, 16'hF71C, 16'hE65A, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hE659, 16'hCD56, 16'hF6DC, 16'hEE9C, 16'hEEDC, 16'hF6DC, 16'hEE9B, 16'hEE9C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF69C, 16'hEE5A, 16'h934E, 16'hEE9B, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hF6DD, 16'hE65B, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'h830D, 16'h000, 16'hD5D9, 16'hF71D, 16'hEEDC, 16'hF6DC,
        16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hDDD8, 16'hD556, 16'hE65A, 16'hF6DC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DD, 16'hCD97, 16'h9411, 16'hFF5D, 16'hC556, 16'h4146, 16'h8B8F, 16'hCD15, 16'hD516, 16'hBC93, 16'h51C8, 16'h73CE, 16'hADD6, 16'h9514, 16'h6C10, 16'hA596, 16'hAD96, 16'hAD97, 16'hAD97, 16'hA596, 16'hADD7, 16'h6BCE, 16'hA452, 16'hFF1D, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hBCD4, 16'h834D, 16'hCD97, 16'hCD96, 16'hCD96, 16'hC556, 16'hDE5A, 16'hF6DC, 16'hF71D, 16'hEE9B, 16'hC556, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCDD7, 16'hBD55, 16'hB514, 16'hD5D8, 16'hD5D7, 16'hDE18, 16'h9410, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h8C10, 16'hCE18, 16'hEEDB, 16'hDE5A, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hDE19, 16'hCD97, 16'hF6DC, 16'hEE9C, 16'hEEDC, 16'hF6DC, 16'hE65B, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC,
        16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hE65A, 16'h82CC, 16'hEE9B, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF6DC, 16'hEE9C, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hE65A, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'h834E, 16'h000, 16'hBD14, 16'hFF1D, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hD597, 16'hCD14, 16'hE61A, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hD5D8, 16'h8B8F, 16'hF6DC, 16'hFF1D, 16'hEE5A, 16'h4A08, 16'h0C3, 16'h3186, 16'h3207, 16'h8491, 16'hA596, 16'hA595, 16'h9D55, 16'h7C92, 16'hA596, 16'hA596, 16'hA596, 16'hA596, 16'hA556, 16'hA596, 16'h94D3,
        16'h7B4E, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hCD97, 16'h6A8A, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hF71C, 16'hD5D8, 16'hC555, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD97, 16'hCD96, 16'hA451, 16'hCDD7, 16'hD5D8, 16'hD618, 16'hC596, 16'h738E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h7B8E, 16'hF71C, 16'hE65A, 16'hE65A, 16'hF71D, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hF6DD, 16'hDDD8, 16'hD5D8, 16'hF6DC, 16'hEE9C, 16'hEEDC, 16'hF6DC, 16'hE65A, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE1A, 16'h6A4A, 16'hE65A, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9B, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hE65A, 16'hEE5B,
        16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hEE9C, 16'hF69C, 16'h8B4E, 16'h58C3, 16'h9BD0, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hD597, 16'hB451, 16'hE619, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hE65A, 16'h838E, 16'hEE9C, 16'hF6DC, 16'hF71D, 16'h838F, 16'h8450, 16'h9D13, 16'h9D54, 16'hAD96, 16'hA555, 16'hA555, 16'h9D55, 16'h4289, 16'h7C50, 16'hAD96, 16'hADD7, 16'hA596, 16'hA596, 16'hADD7, 16'h7C51, 16'h9410, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hDE19, 16'h6A8A, 16'hBD14, 16'hCD97, 16'hC556, 16'hCD97, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71C, 16'hEE9B, 16'hC556, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hD5D7, 16'h9C11, 16'hBD15, 16'hD618, 16'hCDD7, 16'hDE19, 16'h7B4D, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h9C92, 16'hF71D, 16'hD5D8, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hF6DD, 16'hDDD8, 16'hDE19, 16'hF6DC, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hDE19, 16'hE65A,
        16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hE61A, 16'h5186, 16'hDE19, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE5B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hE61A, 16'hE65A, 16'hF6DC, 16'hEE9C, 16'hF69C, 16'hEE9C, 16'hEE9C, 16'hF69C, 16'h834E, 16'h92CC, 16'h82CC, 16'hEE9B, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hD597, 16'hA3CF, 16'hDDD8, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF69C, 16'hEE9B, 16'h834E, 16'hE65B, 16'hF6DD, 16'hF71D, 16'h9C92, 16'h8491, 16'hADD7, 16'hA595,
        16'hA555, 16'hA555, 16'hAD96, 16'h634D, 16'h9C51, 16'h9C51, 16'h4A8A, 16'h8492, 16'h9514, 16'h9D55, 16'h7C11, 16'h3986, 16'hDE59, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hEE9B, 16'h830C, 16'hAC92, 16'hD597, 16'hC556, 16'hD5D8, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hCDD7, 16'hC556, 16'hCD96, 16'hCD96, 16'hCD97, 16'hCD96, 16'hD5D7, 16'hACD3, 16'h93D0, 16'hDE18, 16'hD5D8, 16'hDE59, 16'hAC92, 16'h9CD2, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h8C51, 16'hCE18, 16'hEEDC, 16'hD5D8, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hD5D8, 16'hE65A, 16'hF6DC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hDDD8, 16'hE65A, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE9C, 16'hDDD9, 16'h2000, 16'hD5D8, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hE65B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC,
        16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hE619, 16'hE65A, 16'hF6DC, 16'hEE9C, 16'hF69C, 16'hF69C, 16'hEE9C, 16'hF6DC, 16'h834D, 16'hAB8F, 16'h930D, 16'hD618, 16'hF6DD, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hF6DC, 16'hDDD7, 16'h934D, 16'hD597, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hF69B, 16'h8B8F, 16'hDE19, 16'hF6DD, 16'hFF1D, 16'hC556, 16'h6B8E, 16'hB5D7, 16'hA595, 16'hA596, 16'hADD6, 16'h7C0F, 16'h730C, 16'hEEDC, 16'hFF1D, 16'hCDD8, 16'h9410, 16'h6B0C, 16'h62CB, 16'h838F, 16'hDE59, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF6DC, 16'h938F, 16'h9BD0, 16'hD5D7, 16'hC556, 16'hD5D8, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hE65A, 16'hC556, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD97, 16'hC556, 16'h730C, 16'hCDD7, 16'hD619, 16'hE659, 16'hD618, 16'h6B0C, 16'hF79E, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h7B8E, 16'hEEDB, 16'hE65A, 16'hDDD8, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC,
        16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hD5D8, 16'hEE5B, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hD5D8, 16'hE619, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE9C, 16'hDDD8, 16'h000, 16'hCD97, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hE65A, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hE619, 16'hE619, 16'hEEDC, 16'hEE9C, 16'hF69C, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'h8B8E, 16'hB3D1, 16'hAB8F, 16'hBD15, 16'hF71D, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hDD97, 16'h828B, 16'hCD56, 16'hEE9B, 16'hEE9C,
        16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hF6DC, 16'h93D0, 16'hD5D8, 16'hFF1D, 16'hF6DD, 16'hE69B, 16'h524A, 16'h8C91, 16'hAD95, 16'h9D14, 16'h634D, 16'h730C, 16'hEEDB, 16'hF71D, 16'hF6DC, 16'hFF1D, 16'hFF1D, 16'hEEDC, 16'hEE9C, 16'hFF1D, 16'hF71D, 16'hF6DC, 16'hF71C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hB493, 16'h834D, 16'hCD97, 16'hC556, 16'hD5D8, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF6DC, 16'hCD97, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hD5D7, 16'h838E, 16'hACD3, 16'hDE5A, 16'hE65A, 16'hEE9B, 16'h838E, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8C10, 16'hF71D, 16'hDE19, 16'hE619, 16'hF71D, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hDDD8, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hD597, 16'hE619, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hF69C, 16'hCD97, 16'h000, 16'hCD96, 16'hF6DC, 16'hEE9C, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC,
        16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hE65A, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hF6DC, 16'hDDD8, 16'hDDD8, 16'hF69C, 16'hEE9C, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'h834E, 16'hBC11, 16'hC452, 16'h9C11, 16'hF6DD, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hDD98, 16'h7209, 16'hC514, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hF6DC, 16'h9C11, 16'hC597, 16'hFF1D, 16'hF6DC, 16'hFF1D, 16'hDE5A, 16'h730C, 16'h4A48, 16'h6B0C, 16'hACD4, 16'hEEDC, 16'hF71D, 16'hF6DC, 16'hF6DD, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hFF1D, 16'hCD56, 16'h6A8A, 16'hCD96, 16'hC556, 16'hD5D8, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71C, 16'hDE18, 16'hCD96, 16'hCD96,
        16'hCD96, 16'hCD96, 16'hCD96, 16'hD5D8, 16'hA492, 16'h7B4D, 16'hE65A, 16'hE69B, 16'hEEDC, 16'hB515, 16'h9452, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9C92, 16'hC596, 16'hF71C,
        16'hD5D8, 16'hE69B, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hDE19, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hD597, 16'hDDD9, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hF69C, 16'hCD57, 16'h3800, 16'hBD14, 16'hF6DC, 16'hEE9C, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hE65A, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hF6DC, 16'hD597, 16'hD5D8, 16'hF69C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'h834E, 16'hBC11, 16'hE4D5, 16'h8B4D, 16'hEE9B, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC,
        16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hDDD8, 16'h7208, 16'hB493, 16'hEE5A, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hF6DC, 16'hA452, 16'hBD56, 16'hFF1D, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF6DC, 16'hDE5A, 16'hEEDC, 16'hFF1D, 16'hF71D, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hDE19, 16'h728A, 16'hC555, 16'hCD56, 16'hD5D8, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hEE9B, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD97, 16'hCD97, 16'hCD96, 16'h628A, 16'hD619, 16'hEE9B, 16'hEE9B, 16'hDE59, 16'h6ACB, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h734D, 16'hE69A, 16'hEE9B, 16'hD597, 16'hEE9C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hDE19, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hCD56, 16'hDDD8, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hEEDC, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hF69C, 16'hC516, 16'h5903, 16'hB4D4, 16'hF6DC,
        16'hEE9C, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hE65A, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hD556, 16'hCD56, 16'hF6DC, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF69B, 16'h834D, 16'hBC11, 16'hED56, 16'h930D, 16'hD5D8, 16'hF6DC, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEEDC, 16'hE5D8, 16'h7208, 16'h938F, 16'hE619, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hF6DC, 16'hB493, 16'hB515, 16'hFF1D, 16'hF6DC, 16'hF71D, 16'hF6DC, 16'hF6DD, 16'hF71D, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71C, 16'hEE5A, 16'h72CB,
        16'hB4D3, 16'hCD56, 16'hD5D8, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF6DC, 16'hD5D7, 16'hCD96, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hD5D8, 16'h838E, 16'hBD55, 16'hEEDC, 16'hE69B, 16'hF6DC, 16'h8BCF, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h838F, 16'hEEDC, 16'hE65A, 16'hD5D8, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9B, 16'hDDD8, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hC515, 16'hDDD8, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hF69C, 16'hBCD5, 16'h82CA, 16'hA411, 16'hF6DC, 16'hEE9C, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hE65A, 16'hEE9B, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hCD15, 16'hC514, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hF69B, 16'h7B0C, 16'hBC12,
        16'hED57, 16'hB3D0, 16'hB4D3, 16'hF6DD, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hF6DC, 16'hDDD8, 16'h69C8, 16'h7A8B, 16'hE619, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hBCD4, 16'hACD4, 16'hFF1D, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF69B, 16'h8B4D, 16'hAC51, 16'hCD56, 16'hD5D8, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hDE19, 16'hC596, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hD5D7, 16'hAC93, 16'h838F, 16'hEE9B, 16'hE69B, 16'hF6DC, 16'hC596, 16'h8C51, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB555, 16'hACD3, 16'hF71D, 16'hDDD8, 16'hDE19, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hEE9B, 16'hDDD9, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hC4D4, 16'hDDD8, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC,
        16'hEEDC, 16'hEEDC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hF69C, 16'hAC93, 16'h930C, 16'hA3D0, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hE65A, 16'hEE9B, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hC4D4, 16'hAC52, 16'hF6DC, 16'hEE9B, 16'hF69C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'h7B0C, 16'hCC93, 16'hED57, 16'hCC94, 16'h938E, 16'hF69C, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEEDC, 16'hDD97, 16'h7A8A, 16'h7A49, 16'hDD97, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hC556, 16'hAC93, 16'hFF1D, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC,
        16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'h9BD0, 16'h93CF, 16'hCD56, 16'hD5D8, 16'hF71C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hE69B, 16'hCD96, 16'hCD96, 16'hCD97, 16'hCD97, 16'hCD97, 16'hD597, 16'hC556, 16'h5A49, 16'hDE59, 16'hEEDC, 16'hEE9B, 16'hE69B, 16'h730C, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h8C11, 16'hCDD8, 16'hF6DC, 16'hD5D8, 16'hE65A, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hEE9B, 16'hDDD8, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hBCD4, 16'hD597, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hF69C, 16'hA452, 16'hA38F, 16'h934E, 16'hEE5B, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hE65A, 16'hEE5B, 16'hF6DC, 16'hEE9C, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hEE9C,
        16'hEE9C, 16'hF6DC, 16'hC493, 16'h9BD0, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE5B, 16'h7ACB, 16'hDD16, 16'hED98, 16'hE515, 16'h8B0C, 16'hDE19, 16'hF6DC, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEEDC, 16'hDD97, 16'h828B, 16'h8A8B, 16'hC514, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hCD56, 16'h9C11, 16'hFF1D, 16'hF6DC, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hF6DD, 16'hB4D3, 16'h830D, 16'hCD55, 16'hDE18, 16'hF71D, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hCD97, 16'hCD96, 16'hCD97, 16'hCD97, 16'hD597, 16'hCD97, 16'hD5D8, 16'h7B4D, 16'hBD56, 16'hF6DC, 16'hE69B, 16'hF6DC, 16'h9C51, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h734D, 16'hE69B, 16'hEEDB, 16'hD597, 16'hEE9B, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hEE9B, 16'hDDD8, 16'hEE9B, 16'hEE9B, 16'hEE9B,
        16'hEE9B, 16'hEE9B, 16'hB493, 16'hD597, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hF69C, 16'h93D0, 16'hB410, 16'h930D, 16'hE65A, 16'hF6DC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hE65A, 16'hEE5B, 16'hF6DC, 16'hEE9C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hAC11, 16'h9BCF, 16'hF6DC, 16'hF69C, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hEE5A, 16'h82CB, 16'hE557, 16'hEE1A, 16'hE516, 16'hA38E, 16'hBD15, 16'hF6DD, 16'hEE9B, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hF6DC, 16'hD597, 16'h828A, 16'h9B4D, 16'hA410, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hD598, 16'h93CF, 16'hF71D, 16'hF6DC,
        16'hF71D, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hCD56, 16'h830C, 16'hC515, 16'hDE19, 16'hF71C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hD5D8, 16'hCD96, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hD5D8, 16'hAC93, 16'h83CF, 16'hEEDC, 16'hE69B, 16'hF6DC, 16'hCDD7, 16'h8C51, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8BCF, 16'hF6DC, 16'hE69B, 16'hD597, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hEE5A, 16'hD597, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hAC52, 16'hD556, 16'hEE9B, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'h834E, 16'hCC93, 16'h9B4E, 16'hD5D8, 16'hF6DD, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hE65B, 16'hE65A, 16'hF6DC,
        16'hEE9C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF69C, 16'hF6DC, 16'hAC10, 16'h728B, 16'hC515, 16'hB493, 16'hC516, 16'hC556, 16'hD5D8, 16'hDDD8, 16'h82CB, 16'hEDD8, 16'hFEDD, 16'hE557, 16'hCC93, 16'h9410, 16'hF6DC, 16'hEE9B, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hE5D8, 16'h828A, 16'hBC52, 16'h934E, 16'hE65A, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hDDD8, 16'h938F, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hD5D8, 16'h728A, 16'hBCD4, 16'hDE19, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hE65A, 16'hCD96, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD97, 16'hD5D7, 16'hCD96, 16'h62CB,
        16'hDE5A, 16'hEEDC, 16'hEE9B, 16'hEE9B, 16'h838E, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB555, 16'hB514, 16'hF6DC, 16'hE61A, 16'hCD97, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC,
        16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hE65A, 16'hD597, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'h9BD0, 16'hC514, 16'hEE9B, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'h830D, 16'hD4D4, 16'hAB8F, 16'hC515, 16'hF6DD, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hEE9B, 16'hE65A, 16'hEEDC, 16'hEE9C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE5B, 16'hE5D8, 16'h7ACB, 16'h4946, 16'hA3CF, 16'hB452, 16'hBC93, 16'hB492, 16'hB492, 16'h9BCF, 16'h69C8, 16'hAC10, 16'hCD97, 16'hCC93, 16'hE4D5, 16'h934D, 16'hE65A, 16'hF6DD, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hDD97,
        16'h828A, 16'hD514, 16'h9B4E, 16'hDDD8, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hDDD9, 16'h8B8F, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hF71D, 16'hE619, 16'h82CC, 16'hB493, 16'hE659, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9B, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCDD7, 16'hCDD7, 16'hCD97, 16'hD5D8, 16'h838E, 16'hBD56, 16'hF6DC, 16'hE69B, 16'hF6DD, 16'hA493, 16'hC617, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h8C10, 16'hCDD8, 16'hF6DC, 16'hD5D8, 16'hCD97, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hDE19, 16'hCD55, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'h938F, 16'hBCD4, 16'hEE9B, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hE65A, 16'h830D, 16'hDCD5, 16'hBC11, 16'hAC93, 16'hFEDD, 16'hF6DC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C,
        16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hEE9B, 16'hE65A, 16'hF6DC, 16'hEE9C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hF69C, 16'hE619, 16'h7249, 16'h6A8A, 16'hBCD3, 16'hAC52, 16'hAC52, 16'hA411, 16'hAC51, 16'h934E, 16'h728A, 16'hB410, 16'hB451, 16'hAC10, 16'hAB8F, 16'h7249, 16'hAC92, 16'hE619, 16'hEE9B, 16'hF6DC, 16'hF6DD, 16'hF6DC, 16'hEEDC, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DB, 16'hDDD7, 16'h7A49, 16'hDD56, 16'hA38F, 16'hBD15, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hE619, 16'h938E, 16'hF6DC, 16'hF71C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hE65B, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DD, 16'hEE5A, 16'h934E, 16'hAC51, 16'hE65A, 16'hF71D, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hEEDC,
        16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hD5D8, 16'hCD97, 16'hCD97, 16'hCDD7, 16'hCDD7, 16'hCD97, 16'hD5D8, 16'hAC93, 16'h8BCF, 16'hF6DC, 16'hEE9B, 16'hF6DC, 16'hD5D8, 16'h8C51, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79D, 16'h7B4D,
        16'hE65A, 16'hF6DC, 16'hBD15, 16'hD5D8, 16'hF71D, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hF71D, 16'hD5D8, 16'hBCD4, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF69C, 16'h834D, 16'hAC52, 16'hEE5B, 16'hEEDC, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF69C, 16'hEE5B, 16'h830D, 16'hDD15, 16'hC453, 16'h9BD0, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hEE9C, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hEE9B, 16'hE65A, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hF6DC, 16'hE619, 16'h92CC, 16'h9B8F, 16'hF6DC, 16'hF6DC, 16'hF69C, 16'hE65A, 16'hDE19, 16'hA411, 16'h8ACC, 16'hB411, 16'hA3CF, 16'hA38E, 16'hA38E, 16'h82CB, 16'h4944, 16'h934D, 16'h9B8E, 16'hAC92,
        16'hCD56, 16'hE619, 16'hF69C, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hF69B, 16'hD556, 16'h7A4A, 16'hE597, 16'hC493, 16'hAC51, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hE61A, 16'h8B4E, 16'hEE9C, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hE65A, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF69B, 16'h9BCF, 16'hA411, 16'hE65A, 16'hF6DD, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hDE19, 16'hCD96, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCD97, 16'hD5D7, 16'hC596, 16'h6ACB, 16'hE65A, 16'hEEDC, 16'hEEDB, 16'hEE9B, 16'h7B8E, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD699, 16'h8BCF, 16'hF6DC, 16'hEEDB, 16'hA452, 16'hDE19, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hF71D, 16'hD5D8, 16'hB492, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'h7B0C, 16'h9BCF, 16'hEE5A, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9B, 16'hF69C, 16'hF6DC, 16'hEE9B, 16'hDDD8, 16'hBCD4,
        16'h51C7, 16'hA38F, 16'hA34E, 16'h49C7, 16'hB4D4, 16'hE65A, 16'hF6DC, 16'hEE9C, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hEEDC, 16'hEE9C, 16'hE65A, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hF6DC, 16'hDD97, 16'h9ACC, 16'hA38F, 16'hEE5B, 16'hF69C, 16'hEE9C, 16'hEE9C, 16'hFEDD, 16'hBCD4, 16'hBC11, 16'hFE9B, 16'hF71D, 16'hD515, 16'hCC93, 16'hC493, 16'h6A8A, 16'h8B0C, 16'h934D, 16'h7A49, 16'h71C7, 16'h82CB, 16'h9BCF, 16'hBD14, 16'hDE19, 16'hEE9B, 16'hF6DC, 16'hF6DD, 16'hEEDC, 16'hEE9C, 16'hEE9B, 16'hCD15, 16'h82CB, 16'hE597, 16'hDD56, 16'h938E, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hE65A, 16'h938E, 16'hEE9B, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hE65A, 16'hEE9B, 16'hF6DC,
        16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hB452, 16'h9BD0, 16'hE65A, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hE69A, 16'hCD97, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D8, 16'h730C, 16'hBD56, 16'hF6DC, 16'hE69B, 16'hF71C, 16'hA452, 16'hC617, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'hB514, 16'hF71C, 16'hE65A, 16'h93D0, 16'hEE9B, 16'hF6DD, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hD5D8, 16'hAC52, 16'hF69C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF69C, 16'h8B4E, 16'h728B, 16'hE65A, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hF6DC, 16'hEE9B, 16'hDE19, 16'hC516, 16'hAC12, 16'h9B8F, 16'h8B4D, 16'h4145, 16'h7A8A, 16'hABCF, 16'h830C, 16'hE65A, 16'hF6DC, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hE65B, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hF6DC, 16'hD556, 16'hA30D, 16'hA38F, 16'hEE9B, 16'hF6DC, 16'hF69C, 16'hEE9C,
        16'hF69C, 16'hA411, 16'hCCD3, 16'hFEDD, 16'hFF9F, 16'hF69B, 16'hED97, 16'hFDD9, 16'hA3D0, 16'hBCD4, 16'hEE5A, 16'hD597, 16'hBCD4, 16'h9BD0, 16'h82CC, 16'h7208, 16'h7186, 16'h8B0C, 16'hB493, 16'hD5D8, 16'hF69B, 16'hFEDD, 16'hF69B, 16'hC4D4, 16'h934D, 16'hE597, 16'hED98, 16'h9B4E, 16'hD5D8, 16'hF6DC, 16'hEE9B, 16'hEE9C, 16'hEE5B, 16'h934E, 16'hEE9B, 16'hF71D, 16'hF6DC, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hDE19, 16'hEE9B, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hC515, 16'hA410, 16'hE65A, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hCD97, 16'hCD97, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hDE18, 16'hA452, 16'h9451, 16'hF6DC, 16'hEE9B, 16'hF6DC, 16'hCDD7, 16'h8C51, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h840F, 16'hCDD8, 16'hF6DC, 16'hD5D8, 16'h93D0, 16'hF6DD, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hDDD8, 16'hA411, 16'hF69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF69C, 16'h938E, 16'h50C3, 16'hDE18, 16'hEEDC, 16'hEE9C, 16'hEEDC,
        16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hF6DD, 16'hEE5B, 16'hCD97, 16'hAC52, 16'h9BCF, 16'h8B0C, 16'h8B0C, 16'h9B8F, 16'hAC52, 16'h6A8A, 16'hD515, 16'hF5D8, 16'hAC11, 16'hDDD8, 16'hF69C, 16'hF69C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hE65B, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hF6DC, 16'hC4D4, 16'hB34E, 16'hA38F, 16'hEE9B, 16'hF6DC, 16'hF69C, 16'hF69C, 16'hF69B, 16'h934D, 16'hDD56, 16'hFF5E, 16'hFF5E, 16'hFF1D, 16'hE597, 16'hED98, 16'hD4D4, 16'hA411, 16'hF6DC, 16'hF69C, 16'hF6DC, 16'hF69C, 16'hEE5A, 16'hD5D8, 16'hB493, 16'h8B4E, 16'h6987, 16'h58C3, 16'h82CC, 16'hB493, 16'hDD97, 16'hC492, 16'hABD0, 16'hEDD8, 16'hF5D8, 16'hB411, 16'hBCD4, 16'hF6DC, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'h938E, 16'hEE5B, 16'hF71D, 16'hF6DC, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D,
        16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hE619, 16'hE65A, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hCD56, 16'hB452, 16'hE65A, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hD5D8, 16'hCD97, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D8, 16'hC556, 16'h730C, 16'hE69B, 16'hEEDC, 16'hEEDB, 16'hEE9B, 16'h734D, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h7B8D, 16'hE69B, 16'hF6DC, 16'hBD15, 16'hAC93, 16'hFF1D, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hD5D8, 16'hA3D0, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'h9B8F, 16'h5000, 16'hC515, 16'hF6DC, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hF6DD, 16'hE65A, 16'hC515, 16'h9B8F, 16'h930C, 16'h934D, 16'h934D, 16'h9BCF, 16'hC4D4, 16'hEE5A, 16'hE65A, 16'h830C, 16'hE597, 16'hF5D9, 16'hABD0, 16'hBCD4, 16'hF69C, 16'hEE9B, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9B, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC,
        16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hAC11, 16'hBBD1, 16'hA38F, 16'hEE5B, 16'hF6DC, 16'hF69C, 16'hF6DC, 16'hEE5A, 16'h92CC, 16'hE5D8, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hEE19, 16'hED57, 16'hED97, 16'h930D, 16'hE619, 16'hF69C, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hF69C, 16'hEE9B, 16'hE619, 16'hCD56, 16'hA3D0, 16'h69C7, 16'h6987, 16'h61C8, 16'h934E, 16'hD515, 16'hE597, 16'hDD15, 16'hA411, 16'hF6DC, 16'hEE9B, 16'hEE9C, 16'hF69B, 16'h9B8E, 16'hE65B, 16'hF71D, 16'hF6DC, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hE619, 16'hE61A, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hDDD8, 16'hAC11, 16'hE619, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hDE19, 16'hCD97, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D8, 16'h6ACB, 16'hCDD8, 16'hEEDC, 16'hEE9B, 16'hF6DC, 16'h9C51, 16'hBE17,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h9410, 16'hEEDB, 16'hEE9B, 16'h9C51, 16'hBD15, 16'hFF1D, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hF71D, 16'hD598,
        16'h9B8F, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF69B, 16'h9BCF, 16'h824A, 16'hA410, 16'hF69B, 16'hEEDC, 16'hF6DD, 16'hEE5B, 16'hBCD4, 16'h8B0C, 16'h7A08, 16'h828B, 16'hA3D0, 16'hC515, 16'hDE19, 16'hEE9B, 16'hF69C, 16'hF69C, 16'hDE19, 16'h830C, 16'hE597, 16'hF5D9, 16'hC493, 16'hA411, 16'hF69C, 16'hEE5B, 16'hF69C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF69B, 16'hA38F, 16'hCC93, 16'hABD0, 16'hEE9B, 16'hF6DC, 16'hF69C, 16'hFEDD, 16'hDDD8, 16'h9B0D, 16'hF69B, 16'hFF5F, 16'hFF5E, 16'hFF9F, 16'hF69C, 16'hE557, 16'hF5D8, 16'hB410, 16'hC4D4, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF69C, 16'hF69C, 16'hF69B, 16'hE61A, 16'hD556, 16'h7A8B, 16'h69C8, 16'h7209, 16'h82CC, 16'h9B8E, 16'h724A, 16'hDE19, 16'hF6DC, 16'hEE9C,
        16'hF69B, 16'h938E, 16'hE65A, 16'hF71D, 16'hF6DC, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hE65A, 16'hDE19, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hE619, 16'hB452, 16'hDDD8, 16'hF6DD, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hE65A, 16'hCD97, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hDE18, 16'h9C10, 16'h9C92, 16'hF6DC, 16'hEE9B, 16'hF6DC, 16'hCDD7, 16'h9451, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD14, 16'hB555, 16'hEEDC, 16'hEE9B, 16'h838E, 16'hCDD8, 16'hFF1D, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hF71D, 16'hDDD8, 16'h9B8F, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF69B, 16'h934E, 16'hAB8F, 16'h82CB, 16'hE61A, 16'hF6DC, 16'hCD97, 16'h8B0D, 16'h6146, 16'h82CC, 16'hB4D3, 16'hDE19, 16'hF69B, 16'hF6DC, 16'hF69C, 16'hEE9B, 16'hEE5B, 16'hEE9C, 16'hDE19, 16'h8B0D, 16'hED98, 16'hEDD8, 16'hD516, 16'h938F, 16'hF65B, 16'hEE5B, 16'hF69C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC,
        16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hEE19, 16'hA34E, 16'hDD56, 16'hAC10, 16'hEE9B, 16'hF6DD, 16'hF69C, 16'hFEDD, 16'hC515, 16'hB3D0, 16'hFEDD, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF5E, 16'hED98, 16'hED98, 16'hD515, 16'h9B8F, 16'hF69C, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hF69C, 16'hF69C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF69C, 16'hEDD8, 16'hA38E, 16'hDD56, 16'hD515, 16'hBC52, 16'hB411, 16'h82CB, 16'hA411, 16'hDDD8, 16'hEE9B, 16'hF69B, 16'h9B8F, 16'hE65A, 16'hFF1D, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hE65A, 16'hDE19, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hEEDC, 16'hF71D, 16'hE65A, 16'hB452, 16'hD597, 16'hF6DD, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9B, 16'hCDD7, 16'hCDD7,
        16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D8, 16'hB514, 16'h62CB, 16'hE69B, 16'hEE9B, 16'hEEDC, 16'hEE9B, 16'h7B4E, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h83CF, 16'hD618, 16'hF6DC, 16'hE65A, 16'h6ACB, 16'hE65A, 16'hF71D, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D,
        16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hF71D, 16'hDDD8, 16'h8B4D, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'h8B0D, 16'hC493, 16'hA3CF, 16'h9C10, 16'hA410, 16'h4800, 16'h7A8B, 16'hBD15, 16'hE65A, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF69C, 16'hDE19, 16'h8B0D, 16'hED98, 16'hED98, 16'hE597, 16'h934E, 16'hEE1A, 16'hEE1A, 16'hEE5B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hE5D9, 16'hAB4E, 16'hED98, 16'hAC10, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hFEDD, 16'hAC11, 16'hCC93, 16'hFF1D, 16'hFF9F, 16'hFF5E, 16'hFF9E, 16'hFF9F, 16'hF65A, 16'hED57, 16'hED98, 16'hA34E, 16'hE619, 16'hF6DC, 16'hEE5A, 16'hEE9B, 16'hF69C, 16'hF69C, 16'hF69C, 16'hEE9C, 16'hEE9C,
        16'hEE9B, 16'hF69C, 16'hD515, 16'hA34E, 16'hED98, 16'hF598, 16'hF5D8, 16'hF5D9, 16'hCCD4, 16'hB492, 16'hF69C, 16'hEE9B, 16'hF69C, 16'h9B4E, 16'hE619, 16'hFF1D, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hEE5A, 16'hDDD8, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hEE9B, 16'hB452, 16'hCD56, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hCDD7, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D8, 16'hC596, 16'h3945, 16'hCDD8, 16'hF6DC, 16'hEE9B, 16'hF6DC, 16'h9410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h7B4D, 16'hEE9B, 16'hEEDC, 16'hD5D8, 16'h6ACC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hF71D, 16'hE619, 16'h8B0D, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'h938E, 16'hABD0, 16'h934E, 16'h000, 16'h728A, 16'hBD15, 16'hEE5A, 16'hF6DC, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF69C, 16'hDE19, 16'h8B0D, 16'hED98, 16'hED98, 16'hEDD8, 16'h934E, 16'hDD98, 16'hF65B, 16'hDD97,
        16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hFEDD, 16'hDD97, 16'hB38F, 16'hEDD8, 16'hABD0, 16'hF69B, 16'hF6DC, 16'hF6DC, 16'hF69C, 16'hA34D, 16'hE596, 16'hFF1E, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF1D, 16'hED97, 16'hF5D9, 16'hC412, 16'hBC93, 16'hFEDD, 16'hEE5B, 16'hEE9B, 16'hF69C, 16'hF69C, 16'hF69C, 16'hF69C, 16'hF69C, 16'hEE9B, 16'hFE9C, 16'hBC52, 16'hB3CF, 16'hF61A, 16'hEE1A, 16'hE597, 16'hED98, 16'hE556, 16'hA3D0, 16'hF69B, 16'hEEDC, 16'hF69B, 16'h9B4E, 16'hDE19, 16'hFF1D, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hEE5B, 16'hDDD8, 16'hEEDC, 16'hEE9B, 16'hEEDC, 16'hF6DC, 16'hF71C, 16'hEE9B, 16'hA3D0, 16'hCD15, 16'hEEDC,
        16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hD618, 16'hCD97, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D8, 16'h5A49, 16'hA4D3, 16'hF6DC, 16'hE69B, 16'hF6DC, 16'hBD55, 16'h9C92, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hCE59, 16'h93D0, 16'hF6DC, 16'hEEDC, 16'hBD55, 16'h730D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hF71D, 16'hE61A, 16'h930D, 16'hE65A, 16'hEE9B, 16'hEE9C, 16'hF6DC, 16'hDE18, 16'h59C7, 16'h48C4, 16'h82CB, 16'h6208, 16'hDE19, 16'hFEDC, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF69C, 16'hDDD9, 16'h930D, 16'hEDD8, 16'hED98, 16'hF5D9, 16'hC452, 16'hCD15, 16'hFE9C, 16'hB452, 16'hEE5A, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hFF1D, 16'hCD15, 16'hBC11, 16'hEDD9, 16'hAC10, 16'hF69C, 16'hF6DC, 16'hF6DD, 16'hE61A, 16'hAB8E, 16'hF619, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hEE1A, 16'hED97, 16'hE557, 16'h9B4E, 16'hF69B, 16'hF69C, 16'hE619, 16'hF69B, 16'hF69C, 16'hF69C, 16'hF69C, 16'hF69C, 16'hF69C, 16'hF69B, 16'hA38E, 16'hCC92, 16'hFEDD, 16'hF6DD, 16'hE597, 16'hED98, 16'hF5D8, 16'hA390, 16'hDE19, 16'hF6DC, 16'hF69B, 16'h9B4E, 16'hDDD8, 16'hFF1D, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hEE9B, 16'hDDD8, 16'hEE9B, 16'hEE9B, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF69B, 16'h9BD0, 16'hC4D4, 16'hEE9B, 16'hF71C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71C, 16'hDE19, 16'hCD97, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hCDD7, 16'hDE18, 16'h838E, 16'h6B0C, 16'hEEDC, 16'hEE9B, 16'hEEDC, 16'hE65A, 16'h734D, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'hB514, 16'hF71C, 16'hF6DC, 16'hA492, 16'h9C51, 16'hFF1D, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF6DC, 16'hF71D, 16'hEE5B, 16'h8ACC, 16'hDE59, 16'hFF1D, 16'hE65A, 16'hB493, 16'h6A08, 16'h3000, 16'hABD0, 16'hE557, 16'hA3D0, 16'hBD15, 16'hF69C, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hF69B, 16'hF69B,
        16'hEE9B, 16'hEE9B, 16'hF69C, 16'hE5D8, 16'h930D, 16'hF619, 16'hE598, 16'hEDD8, 16'hDD15, 16'hB412, 16'hFE9D, 16'hBC93, 16'hCD15, 16'hFEDD, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hFEDD, 16'hBC93, 16'hCC93, 16'hEDD9, 16'hB411, 16'hF6DC, 16'hF6DC, 16'hFF1D, 16'hCD56, 16'hB3CF, 16'hF69B, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF1D, 16'hED97, 16'hF5D9, 16'hABD0, 16'hCD56, 16'hFEDD, 16'hDDD8, 16'hEE9B, 16'hF6DC, 16'hF69C, 16'hF69C, 16'hF69C, 16'hF6DC, 16'hEE19, 16'h92CC, 16'hE596, 16'hFF5E, 16'hFF5E, 16'hEDD8, 16'hED98, 16'hF5D9, 16'hBC52, 16'hC515, 16'hF6DC, 16'hF6DB, 16'h9B4E, 16'hD5D8, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D,
        16'hF71D, 16'hEE9B, 16'hDDD8, 16'hEE9B, 16'hEE9B, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'h9BD0, 16'hBC52, 16'hE65A, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hE69B, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hE65A, 16'hCD97, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hDE18, 16'hA492, 16'h000, 16'hDE59, 16'hEEDC, 16'hE69B, 16'hF71C, 16'h8BD0, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h8410, 16'hD619, 16'hEEDC, 16'hF6DC, 16'h838F, 16'hB514, 16'hFF1D, 16'hEEDC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF6DC, 16'hF71D, 16'hEE5B, 16'h930D, 16'hCD97, 16'hC556, 16'h7B0C, 16'h8B8F, 16'hC556, 16'h8B0C, 16'hDD16, 16'hF598, 16'hCCD4, 16'h8B4E, 16'hEE9B, 16'hEE9C, 16'hF69C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hF69B, 16'hF69C, 16'hEE5B, 16'hEE5B, 16'hFEDC, 16'hE5D8, 16'h9B0D, 16'hFEDC, 16'hE5D9, 16'hED98, 16'hED97, 16'hB3D0, 16'hF65B, 16'hDD98, 16'h92CB, 16'hF69B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hF6DD, 16'hF69C, 16'hABD0, 16'hDD15, 16'hF619, 16'hBC52,
        16'hF6DC, 16'hF6DC, 16'hFEDD, 16'hB452, 16'hD493, 16'hFEDD, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF69B, 16'hED98, 16'hD516, 16'h934E, 16'hFEDC, 16'hDDD8, 16'hEE1A, 16'hF6DC, 16'hF69C, 16'hF69C, 16'hF69C, 16'hFEDC, 16'hD515, 16'hA34D, 16'hF65A, 16'hFF5E, 16'hFF5F, 16'hEE5A, 16'hE557, 16'hF5D8, 16'hDD15, 16'hAC11, 16'hF6DC, 16'hF69B, 16'h9B4E, 16'hDE19, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hDDD8, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'h9BD0, 16'hB451, 16'hDE19, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hEE9B, 16'hCD97, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D8, 16'hBD15, 16'h000, 16'hAD14, 16'hEEDC, 16'hE69B, 16'hF71C, 16'hBD55, 16'hA4D3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h7B8E, 16'hEE9B, 16'hEEDC, 16'hEEDB, 16'h6ACB, 16'hC596, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hF6DD, 16'hF69C, 16'hA3CF, 16'h8B8E, 16'hBD15, 16'hDE19, 16'hF6DC, 16'hEE9B, 16'h8B0C, 16'hDD16,
        16'hED57, 16'hED98, 16'h92CC, 16'hDDD8, 16'hF6DC, 16'hEE9C, 16'hF69C, 16'hF69C, 16'hEE9B, 16'hEE5B, 16'hF69B, 16'hF69C, 16'hEE5B, 16'hE61A, 16'hFEDD, 16'hDD98, 16'hA34E, 16'hFF5E, 16'hEE5B, 16'hE597, 16'hF5D9, 16'hBC11, 16'hDD98, 16'hF69B, 16'h8208, 16'hD556, 16'hFEDD, 16'hEE9C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hFF1D, 16'hEE5A, 16'hAB90, 16'hE5D8, 16'hEE1A, 16'hBC52, 16'hF6DC, 16'hF6DD, 16'hF69B, 16'hA34E, 16'hE557, 16'hFF1E, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hEDD9, 16'hEDD8, 16'hA38F, 16'hE619, 16'hE5D9, 16'hDDD8, 16'hFEDD, 16'hF6DC, 16'hF6DC, 16'hF69C, 16'hFEDC, 16'hA3D0, 16'hD4D4, 16'hF6DC, 16'hFF9F, 16'hFF5F, 16'hF6DC, 16'hE597, 16'hED98, 16'hED97, 16'hA38F, 16'hE69B, 16'hFEDC, 16'h930D, 16'hD5D8, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D,
        16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hDE18, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hFEDD, 16'h9BD0, 16'hAC10, 16'hDDD8, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71C, 16'hEE9B, 16'hEE9B, 16'hF71C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D8, 16'hC556, 16'h62CB, 16'h83CF, 16'hE69B, 16'hE69B, 16'hEEDC, 16'hDE5A, 16'h7B8E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h9410, 16'hF71C, 16'hEE9B, 16'hE69B, 16'h5208, 16'hD5D8, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hFEDD, 16'hAC11, 16'hB4D3, 16'hFF1D, 16'hEEDC, 16'hEE9C, 16'hE65A, 16'h930D, 16'hE556, 16'hED98, 16'hF598, 16'hC453, 16'hA411, 16'hF6DC, 16'hEE9B, 16'hF69C, 16'hF69C, 16'hF69C, 16'hEE5A, 16'hF69B, 16'hF69C, 16'hEE5B, 16'hDD98, 16'hFEDD, 16'hDD98, 16'hB411, 16'hFF9E, 16'hF6DD, 16'hED97, 16'hF5D9, 16'hD4D4, 16'hC494, 16'hFEDD, 16'hBC51, 16'h92CB, 16'hF69B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD,
        16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hFF1D, 16'hDD97, 16'hBC11, 16'hF61A, 16'hEE1A, 16'hC493, 16'hFEDD, 16'hFF1E, 16'hE5D8, 16'hB38E, 16'hF61A, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF71D, 16'hEDD8, 16'hDD56, 16'hB452, 16'hE5D8, 16'hD597, 16'hFEDD, 16'hF6DC, 16'hF6DC, 16'hFEDD, 16'hE618, 16'h9B0C, 16'hEDD8, 16'hFF1E, 16'hFF5F, 16'hFF5E, 16'hFF1E, 16'hE5D8, 16'hED98, 16'hF5D8, 16'hABD0, 16'hD5D8, 16'hFEDC, 16'h8ACC, 16'hD597, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hE619, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEEDC, 16'hF6DC, 16'hFF1D, 16'hA411, 16'hA3CF, 16'hD556, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hEE9B, 16'hE65B, 16'hF71C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hD5D7, 16'hCD97, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D8, 16'hCDD7, 16'h838E,
        16'h734C, 16'hD619, 16'hEEDC, 16'hE69B, 16'hEEDC, 16'h7B8E, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'hB515, 16'hF71C, 16'hEEDC, 16'hDE5A, 16'h3986, 16'hDE19, 16'hF6DC, 16'hEEDC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D,
        16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hFF1D, 16'hC4D4, 16'h9BD0, 16'hF6DC, 16'hEE9B, 16'hEEDC, 16'hE65A, 16'h934D, 16'hE556, 16'hF61A, 16'hED98, 16'hED97, 16'h8B0D, 16'hE619, 16'hF6DC, 16'hEE9C, 16'hEE9B, 16'hF69C, 16'hE61A, 16'hEE5A, 16'hF69C, 16'hF69B, 16'hD516, 16'hFEDD, 16'hDD97, 16'hBC92, 16'hFF9F, 16'hFF5E, 16'hEDD9, 16'hED98, 16'hED97, 16'hBC11, 16'hFE9C, 16'hDD97, 16'h9209, 16'hC514, 16'hFF1D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hFF1D, 16'hC4D4, 16'hC452, 16'hF69B, 16'hEE5A, 16'hCCD4, 16'hFF1D, 16'hFF1E, 16'hC4D4, 16'hCC52, 16'hF69C, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hEE5A, 16'hEDD8, 16'hC4D4, 16'hB411, 16'hD556, 16'hFEDD, 16'hF6DC, 16'hF69C, 16'hFEDD, 16'hA3CF, 16'hCC93, 16'hF69B, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hEE5A,
        16'hE597, 16'hF5D9, 16'hC453, 16'hC515, 16'hFEDC, 16'h824A, 16'hD5D7, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hF6DC, 16'hFF1D, 16'hA451, 16'h9B8F, 16'hCD15, 16'hEE9B, 16'hF71D, 16'hF6DC, 16'hF71C, 16'hEE9B, 16'hE65A, 16'hF71C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hDE18, 16'hCD96, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D8, 16'hD5D8, 16'h8BD0, 16'h9C92, 16'hBD56, 16'hF71C, 16'hE69B, 16'hF6DC, 16'hACD3, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h8C10, 16'hD618, 16'hF6DC, 16'hF6DC, 16'hD5D8, 16'h3946, 16'hE65A, 16'hF6DC, 16'hEE9B, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hFF1D, 16'hDD57, 16'h82CC, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hE65A, 16'h934D, 16'hE556, 16'hF69C, 16'hF65A, 16'hED98, 16'hC494, 16'hA411, 16'hFEDD, 16'hEE9C, 16'hF69C, 16'hF6DC, 16'hEE5A, 16'hDDD8, 16'hFEDC, 16'hFEDC, 16'hCD15, 16'hF65B, 16'hDD97, 16'hC4D4, 16'hFF9F, 16'hFF9E, 16'hF69B, 16'hED98, 16'hF5D9, 16'hB3D1, 16'hE619, 16'hF65A, 16'hBC11, 16'hAB8F, 16'hE619, 16'hFEDD, 16'hF6DC, 16'hF6DC, 16'hF6DC,
        16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hFEDD, 16'hB451, 16'hD4D5, 16'hFEDC, 16'hE619, 16'hCD15, 16'hFF1E, 16'hF69C, 16'hAB8F, 16'hE556, 16'hFF1D, 16'hFF9F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hEE5A, 16'hF65A, 16'hB411, 16'hC4D4, 16'hFEDD, 16'hF6DC, 16'hFF1D, 16'hCD15, 16'hB3D0, 16'hF5D8, 16'hF6DD, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hF6DD, 16'hED97, 16'hF5D9, 16'hD4D5, 16'hB452, 16'hF69B, 16'h71C8, 16'hD5D7, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hE65A, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hFF1D, 16'hAC93, 16'h8B0D, 16'hCD15, 16'hE65A, 16'hF71D, 16'hF6DC, 16'hF71C, 16'hEE9C, 16'hDE19, 16'hF6DC, 16'hF6DC,
        16'hF6DC, 16'hF6DC, 16'hF71C, 16'hDE19, 16'hCD96, 16'hCDD7, 16'hD5D7, 16'hD5D7, 16'hD5D8, 16'hD5D8, 16'hDE18, 16'h9410, 16'hAD15, 16'hA493, 16'hEEDC, 16'hE69B, 16'hEEDC, 16'hD619, 16'h8410, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h838E, 16'hEEDB, 16'hEE9B, 16'hF71C, 16'hC597, 16'h3946, 16'hE65B, 16'hF6DC, 16'hEE9B,
        16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hFF1D, 16'hE5D9, 16'h6986, 16'hDE19, 16'hF6DC, 16'hF6DC, 16'hE65A, 16'h9B4E, 16'hE557, 16'hF69C, 16'hFF5E, 16'hE557, 16'hEDD8, 16'h9B4E, 16'hDDD9, 16'hF6DD, 16'hF69C, 16'hF69C, 16'hF69B, 16'hD515, 16'hF69B, 16'hFF1D, 16'hD556, 16'hE619, 16'hDD98, 16'hCD56, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hEDD9, 16'hF5D9, 16'hD4D4, 16'hC4D5, 16'hFEDD, 16'hC493, 16'hC411, 16'hBC11, 16'hFEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF6DD, 16'hFF1D, 16'hF69B, 16'hB3D0, 16'hE557, 16'hFF1D, 16'hDDD8, 16'hD556, 16'hFF5F, 16'hDD98, 16'hB3CF, 16'hEE19, 16'hFF5E, 16'hFF9F, 16'hFF5D, 16'hEE9B, 16'hE619, 16'hDDD8, 16'hD596, 16'hD556, 16'hCD56, 16'hC515, 16'hD597, 16'hDE1A, 16'hE65A, 16'hEDD8, 16'hBC52, 16'hCD15,
        16'hFF1E, 16'hFEDD, 16'hD556, 16'hABCF, 16'hED97, 16'hEE1A, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hEDD9, 16'hEDD8, 16'hE556, 16'hB451, 16'hF65A, 16'h7187, 16'hD597, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hE65A, 16'hE65B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hFF1D, 16'hB4D4, 16'h7ACC, 16'hCD15, 16'hDDD8, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hDE19, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hE65A, 16'hCD96, 16'hCDD7, 16'hD5D7, 16'hD5D8, 16'hD5D8, 16'hD5D7, 16'hDE19, 16'h9C51, 16'hB596, 16'hA4D3, 16'hDE59, 16'hEEDC, 16'hE69B, 16'hEEDB, 16'h7B8E, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h9C51, 16'hF71C, 16'hE69B, 16'hF71C, 16'hB514, 16'h628A, 16'hF6DC, 16'hEE9C, 16'hEE9B, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hEE5A, 16'h6905, 16'hC515, 16'hF71D, 16'hF6DC, 16'hE65A, 16'h9B4E, 16'hED57, 16'hF69B, 16'hFF9F, 16'hEE1A, 16'hED97, 16'hDD56, 16'h9BCF, 16'hF69C, 16'hF69C, 16'hF69C, 16'hFEDD, 16'hCCD5, 16'hDDD8, 16'hFF1D, 16'hE5D9, 16'hDD97, 16'hDD98, 16'hD597, 16'hFFDF, 16'hFF9F, 16'hFF9F,
        16'hF6DC, 16'hED98, 16'hED97, 16'hBC11, 16'hFE9C, 16'hDD97, 16'hC452, 16'hC452, 16'hD556, 16'hFF1D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF6DD, 16'hFF1E, 16'hE619, 16'hB38F, 16'hF5D9, 16'hFF5E, 16'hD556, 16'hE5D8, 16'hFF1E, 16'hBC11, 16'hD4D4, 16'hF69B, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hF71D, 16'hF6DC, 16'hEE9C, 16'hE65A, 16'hDE19, 16'hCDD8, 16'hBCD4, 16'h934E, 16'hAC11, 16'hC4D4, 16'hA34E, 16'hAB4E, 16'hEDD9, 16'hFE9B, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5F, 16'hF65B, 16'hED98, 16'hED57, 16'hBC11, 16'hEE19, 16'h7105, 16'hD597, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF6DC,
        16'hFF1D, 16'hBD15, 16'h7A8B, 16'hCD15, 16'hD597, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hDE19, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hEE9B, 16'hCD96, 16'hCD97, 16'hCD97, 16'hD5D7, 16'hD5D8, 16'hD5D8, 16'hDE18, 16'hACD3, 16'hA514, 16'hAD15, 16'hC5D7, 16'hF6DC, 16'hE69B, 16'hF71C, 16'h9C92, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hB555, 16'hB515, 16'hF71D, 16'hEE9B, 16'hF71C, 16'h9C92, 16'h730C, 16'hF6DC, 16'hEE9B, 16'hE65B, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF71D, 16'hF69B, 16'h8A8A, 16'h938E, 16'hF6DC, 16'hF71C, 16'hDE19, 16'h9B8E, 16'hED98, 16'hF69B, 16'hFFDF, 16'hFF5E, 16'hE597, 16'hF619, 16'hBC93, 16'hB492, 16'hFEDD, 16'hF69C, 16'hFEDC, 16'hE5D9, 16'hBC92, 16'hFF1D, 16'hF69B, 16'hDD97, 16'hD557, 16'hDDD8, 16'hFF9F, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hEDD8, 16'hF5D8, 16'hCC93, 16'hDD97, 16'hFEDC, 16'hB411, 16'hE556, 16'hA38E, 16'hEE5B, 16'hFEDD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF69C, 16'hFEDD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF6DD, 16'hFF1E, 16'hD556, 16'hC411, 16'hF65A, 16'hFF9F, 16'hC493, 16'hEE5A, 16'hEE1A, 16'hB38F, 16'hEDD8, 16'hF71D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1D, 16'hEE5A, 16'hE619, 16'hDDD8, 16'hCD56, 16'hCCD5, 16'hDDD8, 16'hF6DC, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hF6DC, 16'hEDD8, 16'hED98, 16'hC493, 16'hE597, 16'h6800, 16'hDD97, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hE65A, 16'hEE5A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hFF1D, 16'hC556, 16'h6208, 16'hCCD5, 16'hCD15, 16'hF6DC, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hDE19, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9B, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCDD7, 16'hD5D8, 16'hD5D8, 16'hD618, 16'hC555, 16'h8C10, 16'hC5D8, 16'hA4D3, 16'hF71C, 16'hE69B, 16'hEEDC, 16'hBD56, 16'h9C92, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h8C10, 16'hD618, 16'hF71C, 16'hEEDB, 16'hF71C, 16'h83CF, 16'h7B4E, 16'hF6DC, 16'hEE5B, 16'hE65A, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFEDC, 16'hA38F, 16'h6146, 16'hE65A, 16'hFF1D, 16'hDDD8, 16'hA38F, 16'hED98, 16'hF6DC, 16'hFFDF, 16'hFF9F, 16'hF6DC, 16'hED98, 16'hF619, 16'hABD1, 16'hBCD4,
        16'hFE9C, 16'hFEDD, 16'hFEDD, 16'hB452, 16'hF69B, 16'hF69A, 16'hBC52, 16'hB411, 16'hC493, 16'hE5D8, 16'hDDD9, 16'hEE5B, 16'hF6DC, 16'hFEDC, 16'hEE19, 16'hE597, 16'hC453, 16'hFF1D, 16'hD556, 16'hD4D4, 16'hE556, 16'hB411, 16'hFEDD, 16'hF6DD, 16'hF6DC, 16'hF6DD, 16'hEE9B, 16'hF6DD, 16'hFF1D, 16'hFEDD, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF6DD, 16'hFEDD, 16'hBC93, 16'hDD15, 16'hF6DC, 16'hFF5E, 16'hC493, 16'hFE9C, 16'hC493, 16'hD4D4, 16'hF619, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF1D, 16'hEE5A, 16'hDD97, 16'hBCD3, 16'hB411, 16'hA3D0, 16'h8B0D, 16'h6A49, 16'h7ACC, 16'h8B4E, 16'h9BCF, 16'hB4D4, 16'hDE5A, 16'hF71D, 16'hFF5E, 16'hF71D, 16'hF6DC, 16'hF71D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hEDD9, 16'hED98, 16'hD4D4, 16'hD516, 16'h7000, 16'hD556, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D,
        16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hEE5B, 16'hE65A, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hFF1D, 16'hCD96, 16'h61C8, 16'hCCD5, 16'hC515, 16'hEE5B, 16'hF71D, 16'hF6DC, 16'hF6DD, 16'hDE19, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hCD97, 16'hCD96, 16'hCD97, 16'hCD97, 16'hD5D8, 16'hD5D8, 16'hD618, 16'hD5D7, 16'h7B8E, 16'hD69A, 16'h9451, 16'hEEDB, 16'hEEDB, 16'hEEDC, 16'hDE5A, 16'h7B8E, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'h7B8E, 16'hEEDB, 16'hEEDC, 16'hEEDC, 16'hEEDB, 16'h5249, 16'h83CF, 16'hF6DC, 16'hE65A, 16'hE61A, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hFF1D, 16'hBC52, 16'h4800, 16'hD597, 16'hFF5E, 16'hD596, 16'hABD0, 16'hED98, 16'hF6DC, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hEE1A, 16'hE598, 16'hEDD9, 16'hB411, 16'hA38F, 16'hCD15, 16'hEE5A, 16'hBC52, 16'h9B0D, 16'hBC93, 16'hC556, 16'hE65A, 16'hF71D, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF71C, 16'hF619, 16'hC493, 16'hE61A, 16'hFF1D, 16'hBC12, 16'hFE19, 16'hCC52, 16'hBC94, 16'hFF1D, 16'hF6DC, 16'hFEDD, 16'hF69C, 16'hF69C, 16'hFF1D, 16'hF6DC, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFEDD, 16'hFF1D, 16'hF69C, 16'hEE19, 16'hBC51, 16'hED97,
        16'hFF1D, 16'hF71D, 16'hD4D5, 16'hEE1A, 16'hB38F, 16'hF597, 16'hF69B, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hEE5A, 16'hD515, 16'hAB4E, 16'h7186, 16'h58C3, 16'h4882, 16'h3000, 16'h2800, 16'h000, 16'h000, 16'h1000, 16'h800, 16'h000, 16'h000, 16'h1800, 16'h83CF, 16'hB596, 16'hDEDB, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hFF5E, 16'hFF9F, 16'hF71D, 16'hEE19, 16'hED97, 16'hD4D4, 16'hC493, 16'h9A4B, 16'hD556, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hEE9B, 16'hE65A, 16'hE65B, 16'hEE9B, 16'hEE9B, 16'hEEDC, 16'hFF1D, 16'hCD97, 16'h5986, 16'hC4D4, 16'hC515, 16'hE619, 16'hF71D, 16'hF6DC, 16'hF6DD, 16'hE61A, 16'hE65A, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hD5D7, 16'hCD96, 16'hCD97, 16'hCD97, 16'hD5D7, 16'hD5D8, 16'hD5D8, 16'hDE19, 16'h8BCF, 16'hD69A, 16'h9C92, 16'hDE59, 16'hEEDC, 16'hE69B, 16'hEEDC, 16'h83CF,
        16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h9410, 16'hF71D, 16'hEEDC, 16'hF6DC, 16'hE69A, 16'h000, 16'h9410, 16'hF6DC, 16'hE619, 16'hE619, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hFF1D, 16'hCD15, 16'h5800, 16'hB452,
        16'hFF5E, 16'hC515, 16'hBC11, 16'hF5D9, 16'hFF1D, 16'hFFDF, 16'hFF9F, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hF61A, 16'hE598, 16'hA34E, 16'hA38F, 16'hB493, 16'hDDD9, 16'hF6DD, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9F, 16'hF6DC, 16'hE597, 16'hC453, 16'hFF5E, 16'hD556, 16'hDD56, 16'hFE59, 16'hBBD0, 16'hCD15, 16'hFF1D, 16'hF6DC, 16'hFEDD, 16'hEE5A, 16'hFF1D, 16'hF69B, 16'hF6DC, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hE5D8, 16'hDD97, 16'hD4D4, 16'hEDD9, 16'hFF5F, 16'hEE9B, 16'hDD16, 16'hCCD4, 16'hD494, 16'hF619, 16'hFF5E, 16'hFF9F, 16'hFF5F, 16'hF71D, 16'hEE9B, 16'hE5D8, 16'hABD0, 16'h6A08, 16'h4945, 16'h4905, 16'h5145, 16'h4945, 16'h5186, 16'h5986, 16'h5146, 16'h4945, 16'h4945, 16'h4945, 16'h4145, 16'h3945, 16'h2882, 16'h000, 16'h000, 16'h000, 16'h6ACB, 16'hC596, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'hDE19, 16'hF6DB, 16'hED97, 16'hD493, 16'hBC11, 16'hB3D0, 16'hD556, 16'hFF5E,
        16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hEE9B, 16'hE65A, 16'hE65B, 16'hEE9B, 16'hEE9B, 16'hEEDC, 16'hFF1D, 16'hD5D7, 16'h5987, 16'hC494, 16'hC4D5, 16'hD5D8, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hE65A, 16'hE65A, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hD5D8, 16'hCD96, 16'hCD97, 16'hCD97, 16'hCDD7, 16'hD618, 16'hD618, 16'hDE59, 16'h9C51, 16'hCE59, 16'hBD96, 16'hBD96, 16'hF71C, 16'hE69B, 16'hF71C, 16'hA4D3, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB595, 16'hB514, 16'hF71D, 16'hEEDB, 16'hF71C, 16'hD5D8, 16'h000, 16'h9411, 16'hF6DC, 16'hDDD8, 16'hE619, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hFF1E, 16'hDD97, 16'h8187, 16'h8A8B, 16'hEE9B, 16'hCD56, 16'hC453, 16'hF619, 16'hFF9E, 16'hFF9F, 16'hF71D, 16'hFF5E, 16'hFF9F, 16'hFF5E, 16'hCD56, 16'hCD56, 16'hF71C, 16'hFF5E, 16'hE69B, 16'hD619, 16'hC556, 16'hAC52, 16'hB410, 16'hB3D0, 16'hBBD1, 16'hC453, 16'hDD97, 16'hF69B, 16'hFF1E, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hF69B, 16'hCC94, 16'hE619, 16'hFEDC, 16'hCC94, 16'hF65A, 16'hF5D8, 16'hB3D0, 16'hD556, 16'hFF1E, 16'hFF1D, 16'hE619, 16'hF69C, 16'hF69B, 16'hE619, 16'hFF1E,
        16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hEE9B, 16'hDD15, 16'hD515, 16'hE597, 16'hEE5A, 16'hFFDF, 16'hE5D8, 16'hDC94, 16'hCC93, 16'hED98, 16'hEE5A, 16'hFF9F, 16'hFF5E, 16'hF71C, 16'hF6DC, 16'hF6DC, 16'hD556, 16'h828A, 16'h6145, 16'h7208, 16'h7208, 16'h69C8, 16'h5145, 16'h4000, 16'h3000, 16'h3801, 16'h4104, 16'h4104, 16'h3904, 16'h3903, 16'h3903, 16'h3904, 16'h3945, 16'h3945, 16'h3104, 16'h000, 16'h000, 16'h51C6, 16'hC555, 16'hBD56, 16'h9BCF, 16'hEEDC, 16'hFF5E, 16'hE557, 16'hA30D, 16'hDD57, 16'hBC11, 16'hCD56, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hEE5B, 16'hE65A, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hF6DC, 16'hFF1D, 16'hDDD8, 16'h5987, 16'hBC53, 16'hCCD5, 16'hCD97, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hE65B, 16'hE619, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hDE18, 16'hCD96, 16'hCD97, 16'hCDD7,
        16'hCD97, 16'hD5D8, 16'hD618, 16'hDE59, 16'hACD3, 16'hBD96, 16'hDEDB, 16'h9C92, 16'hF71C, 16'hEE9B, 16'hF6DC, 16'hCDD7, 16'h9451, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h8C10, 16'hCDD8, 16'hF71D, 16'hEEDB, 16'hF71D, 16'hBD55, 16'h000, 16'hA492, 16'hF6DC, 16'hD557, 16'hE619, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D,
        16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hFF1D, 16'hE619, 16'h8A49, 16'h9A8B, 16'hC515, 16'hDD97, 16'hCC93, 16'hF65A, 16'hFF5E, 16'hF71D, 16'hFF9E, 16'hFF9F, 16'hFF5E, 16'hEE9B, 16'hF6DC, 16'hF71D, 16'hC597, 16'h734D, 16'h1800, 16'h000, 16'h000, 16'h2000, 16'h4800, 16'h58C4, 16'h7146, 16'h9A8B, 16'hAB0D, 16'hC3D1, 16'hE5D8, 16'hEE5B, 16'hF69B, 16'hFF5E, 16'hFF5E, 16'hEE19, 16'hC453, 16'hFF5E, 16'hDD97, 16'hE598, 16'hF65A, 16'hF5D9, 16'hB411, 16'hD597, 16'hFF5F, 16'hEE9B, 16'hDD97, 16'hFF1D, 16'hD4D4, 16'hFEDD, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hDD56, 16'hDD16, 16'hD4D5, 16'hED97, 16'hF6DC, 16'hFF5E, 16'hDD15, 16'hC3D0, 16'hE597, 16'hE5D8, 16'hF71D, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hF6DC, 16'hBC93, 16'h8249, 16'h7A09, 16'h8249, 16'h69C7, 16'h4801, 16'h2800, 16'h4905, 16'h830D, 16'h9BCF, 16'h834D, 16'h6249, 16'h4145, 16'h4945, 16'h4945, 16'h4145, 16'h4104, 16'h3904, 16'h38C3, 16'h30C3, 16'h30C3, 16'h3104,
        16'h2001, 16'h000, 16'h000, 16'hC556, 16'hE659, 16'hD597, 16'hD4D4, 16'hD4D5, 16'hFE5B, 16'hAB8F, 16'hD597, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hF6DC, 16'hF71D, 16'hDE19, 16'h59C7, 16'hBC52, 16'hCCD5, 16'hCD56, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hEE9B, 16'hDE19, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hDE19, 16'hCD96, 16'hCD97, 16'hCDD7, 16'hC596, 16'hCD97, 16'hD618, 16'hDE19, 16'hC596, 16'h9C92, 16'hEF5D, 16'h9411, 16'hEEDC, 16'hEEDB, 16'hEEDC, 16'hE65A, 16'h7B8E, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h7B8E, 16'hE69B, 16'hEEDC, 16'hEEDB, 16'hF71C, 16'hA493, 16'h000, 16'hA493, 16'hF6DC, 16'hCD56, 16'hE65A, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF69B, 16'h8A4A, 16'hBB90, 16'hA38F, 16'hD556, 16'hDD15, 16'hF69B, 16'hFF5E, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hEEDC, 16'hACD4, 16'h2880, 16'h000, 16'h000, 16'h2882, 16'h4145, 16'h4145, 16'h4145, 16'h4104, 16'h4104, 16'h5145, 16'h5945, 16'h69C7, 16'h71C8, 16'hBC51, 16'hEE19, 16'hF6DC, 16'hF6DC, 16'hF71E, 16'hFF1D, 16'hDD16, 16'hD556,
        16'hFF1D, 16'hD556, 16'hFEDC, 16'hF619, 16'hF61A, 16'hBC11, 16'hD556, 16'hFF1D, 16'hD4D5, 16'hF6DC, 16'hC4D4, 16'hCD15, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hF69C, 16'hCCD4, 16'hD556, 16'hDD16, 16'hEDD8, 16'hFF9F, 16'hEE9B, 16'hC38F, 16'hE5D8, 16'hEE5A, 16'hF69B, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hDE19, 16'hA30D, 16'h89C7, 16'h8A8A, 16'h79C8, 16'h3800, 16'h4104, 16'h830D, 16'hAC92, 16'hD596, 16'hCD56, 16'h93CF, 16'h41C7, 16'h3145, 16'h2103, 16'h20C3, 16'h2903, 16'h3104, 16'h3103, 16'h30C3, 16'h3904, 16'h4104, 16'h4104, 16'h30C3, 16'h28C3, 16'h2904, 16'h18C3, 16'h801, 16'h9411, 16'hB4D3, 16'hCD14, 16'hEDD9, 16'hFE5B, 16'hAB8F, 16'hD597, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hF6DC, 16'hF71D, 16'hE65A, 16'h59C8, 16'hBC52, 16'hCCD5, 16'hCD15, 16'hE65A, 16'hF71C,
        16'hF6DC, 16'hEE9B, 16'hDE19, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hDE59, 16'hCD96, 16'hCDD7, 16'hCDD7, 16'hC596, 16'hB514, 16'hD618, 16'hD618, 16'hCDD8, 16'h83CF, 16'hF79E, 16'h9451, 16'hDE59, 16'hEEDC, 16'hEE9B, 16'hEEDC, 16'h838E, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8BD0, 16'hF71C, 16'hEEDC, 16'hEEDC, 16'hF71C, 16'h9410, 16'h5A8A,
        16'h9C52, 16'hF69C, 16'hCD15, 16'hE65A, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hA34E, 16'hBB90, 16'hCCD4, 16'hA38F, 16'hE557, 16'hF69B, 16'hFF9F, 16'hEF1C, 16'hEF1C, 16'hFF9E, 16'hBD56, 16'h1000, 16'h000, 16'h1000, 16'h3104, 16'h3104, 16'h4144, 16'h4945, 16'h5145, 16'h5145, 16'h5986, 16'h6186, 16'h6987, 16'h69C7, 16'h71C8, 16'h79C8, 16'h7987, 16'h9B0D, 16'hDD97, 16'hF71D, 16'hFF9F, 16'hFF5E, 16'hF65A, 16'hCC93, 16'hE61A, 16'hF69B, 16'hE619, 16'hFEDC, 16'hEDD8, 16'hF65A, 16'hC452, 16'hBC12, 16'hD4D4, 16'hCCD4, 16'hEE19, 16'hB3D0, 16'hD557, 16'hF6DC, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hCD15, 16'hE5D8, 16'hEE5A, 16'hE598, 16'hF69C, 16'hFF5F, 16'hD516, 16'hE5D8, 16'hFF1D, 16'hEE19, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hEE9B, 16'hCCD4, 16'hAB4E, 16'h9ACC, 16'h7987, 16'h82CB, 16'hA451, 16'hCD55, 16'hD5D7, 16'hE618, 16'hC554, 16'h3104, 16'h000,
        16'h101, 16'h1984, 16'h29C5, 16'h29C5, 16'h2A06, 16'h29C5, 16'h2A06, 16'h21C5, 16'h1943, 16'h2103, 16'h2082, 16'h3904, 16'h3904, 16'h28C3, 16'h28C3, 16'h2082, 16'h000, 16'h3986, 16'h9C10, 16'hB452, 16'hE5D8, 16'hAB8F, 16'hD597, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hE65B, 16'hEE5A, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hF6DC, 16'hF71D, 16'hEE9B, 16'h6249, 16'hB412, 16'hCCD5, 16'hCD55, 16'hDE19, 16'hF6DC, 16'hF71D, 16'hEE9C, 16'hDE19, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hF71D, 16'hDE5A, 16'hCD96, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hA492, 16'hD5D8, 16'hD618, 16'hD618, 16'h7B8E, 16'hF75D, 16'hA514, 16'hCDD7, 16'hEEDC, 16'hE69B, 16'hF6DC, 16'h9C52, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC5D7, 16'hA493, 16'hF71D, 16'hEEDC, 16'hF6DC, 16'hE69B, 16'h838F, 16'hA4D3, 16'h9411, 16'hEE9B, 16'hC4D5, 16'hE65A, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1E, 16'hBC92, 16'hAACD, 16'hEDD8, 16'hB411, 16'hDD56, 16'hF65A, 16'hFF5D, 16'hE69A, 16'h9C51, 16'h62CA, 16'h000, 16'h1841, 16'h2904, 16'h30C3, 16'h4945, 16'h4144, 16'h3000, 16'h38C1, 16'h4986, 16'h4145, 16'h4945, 16'h4144,
        16'h4945, 16'h5186, 16'h61C7, 16'h69C8, 16'h7A49, 16'h8A4A, 16'hB30D, 16'hCC52, 16'hEE5B, 16'hFF5E, 16'hF69B, 16'hF61A, 16'hCC93, 16'hEE59, 16'hE619, 16'hF71D, 16'hF69C, 16'hEDD8, 16'hFE9B, 16'hE619, 16'hCC94, 16'hCCD4, 16'hD515, 16'hE597, 16'hDD98, 16'hBC52, 16'hD515, 16'hDD97, 16'hDD97, 16'hDD97, 16'hE5D9, 16'hF69C, 16'hF65A, 16'hF69B, 16'hFF9F, 16'hFF5E, 16'hFF1D, 16'hFF9F, 16'hF6DC, 16'hFF1D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hE65A, 16'hCCD5, 16'hCCD4, 16'h79C7, 16'hB492, 16'hD5D7, 16'hDE18, 16'hD5D7, 16'hD5D7, 16'hBD14, 16'h000, 16'h902, 16'h3A47, 16'h3A47, 16'h42C9, 16'h4B0A, 16'h534B, 16'h538B, 16'h538B, 16'h534B, 16'h534B, 16'h4B09, 16'h4288, 16'h29C5, 16'h2103, 16'h800, 16'h28C3, 16'h4104, 16'h30C3, 16'h3144, 16'h000, 16'h000, 16'h4146, 16'hAC11, 16'h9B0D, 16'hDE19, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hE65A, 16'hEE5A,
        16'hEE5A, 16'hEE5B, 16'hEE5B, 16'hF6DC, 16'hF6DD, 16'hEE9B, 16'h6A8A, 16'hABD1, 16'hCCD5, 16'hCD56, 16'hD5D8, 16'hF6DC, 16'hF6DD, 16'hEEDC, 16'hDE19, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hE65A, 16'hCD97, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'h9410, 16'hC596, 16'hDE19, 16'hDE59, 16'h83CF, 16'hE6DB, 16'hC618, 16'hACD4, 16'hEEDC, 16'hE69B, 16'hEEDC, 16'hBD55, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'hC596, 16'hF71D, 16'hEEDC, 16'hF71C, 16'hD659, 16'h8C11, 16'hBDD7, 16'h8BD0, 16'hEE5B, 16'hC4D5, 16'hE65A, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1E, 16'hCD56, 16'hA24B, 16'hF65A, 16'hEE9A, 16'hD556, 16'hF619, 16'hF65A, 16'hEE9C, 16'h738E, 16'h000, 16'h2945, 16'h2082, 16'h4145, 16'h4104, 16'h000, 16'h1800, 16'h72CB, 16'h730C, 16'h5A49, 16'h2103, 16'h18C3, 16'h1103, 16'h1943, 16'h1984, 16'h1944, 16'h2144, 16'h20C2, 16'h4145, 16'h82CB, 16'hBB90, 16'hE557, 16'hFF5E, 16'hFF1E, 16'hF69B, 16'hF659, 16'hD515, 16'hD556, 16'hE619, 16'hFF9F, 16'hF6DC, 16'hEE19, 16'hFEDC, 16'hFF5E, 16'hFF5E, 16'hEE9B, 16'hE619, 16'hFF5E, 16'hFF5E, 16'hF71D, 16'hFF5E, 16'hFF5D, 16'hFF5E, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hEE9B, 16'hEE9B,
        16'hFF1D, 16'hB493, 16'hBCD3, 16'hDE18, 16'hD5D7, 16'hD596, 16'hD5D7, 16'hCD96, 16'h4A07, 16'h1103, 16'h4288, 16'h4B0A, 16'h5B8C, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h534B, 16'h4B0A, 16'h3206, 16'h000, 16'h38C3, 16'h4985, 16'h3904, 16'h2882, 16'h28C3, 16'h000, 16'h41C7, 16'h6A08, 16'hE61A, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hE65A, 16'hEE5A, 16'hEE5A, 16'hEE5B, 16'hEE9B, 16'hF6DC, 16'hF6DD, 16'hEE9B, 16'h6249, 16'hAC11, 16'hC4D4, 16'hCD56, 16'hD597, 16'hEEDC, 16'hF71D, 16'hF6DC, 16'hDE19, 16'hEE9B, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hE65A, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D8, 16'h9410, 16'hACD3, 16'hDE59, 16'hDE59, 16'h9451, 16'hCE59, 16'hE71C, 16'h9451, 16'hEEDC, 16'hE69B, 16'hEEDC, 16'hD618, 16'h83CF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h8410, 16'hD619, 16'hF71C, 16'hEEDC, 16'hF71D, 16'hC5D7, 16'hAD15, 16'hCE19, 16'h8BD0, 16'hEE5A, 16'hC515, 16'hEE5A, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hDDD8, 16'h9209, 16'hEDD8, 16'hFF5D, 16'hF69B, 16'hDD56, 16'hD556, 16'h5208, 16'h000, 16'h2904,
        16'h30C2, 16'h4145, 16'h1000, 16'h1800, 16'h8B8E, 16'hBD14, 16'h9410, 16'h4207, 16'h1984, 16'h2205, 16'h2A46, 16'h3247, 16'h3247, 16'h3A87, 16'h3A88, 16'h3A47, 16'h3A06, 16'h1903, 16'h51C7, 16'hB451, 16'hD556, 16'hF6DC, 16'hFF9F, 16'hFF5E, 16'hFF1E, 16'hFF5F, 16'hEE9B, 16'hE619, 16'hFF5E, 16'hFF9F, 16'hFF1E, 16'hF6DC, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hF75E, 16'hDE19, 16'hD596, 16'hD5D6, 16'hD5D7, 16'hD5D7, 16'hDDD7, 16'h93CF, 16'h000, 16'h4AC9, 16'h5B8C, 16'h640D, 16'h63CD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h538C, 16'h3A88, 16'h1102, 16'h28C3, 16'h4986, 16'h4946, 16'h3903, 16'h28C3, 16'h000, 16'h2000, 16'hE65A, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D,
        16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hE65A, 16'hEE5A, 16'hEE5A, 16'hEE5B, 16'hEE9B, 16'hF6DC, 16'hF6DD, 16'hEE9B, 16'h6249, 16'hAC11, 16'hCCD4, 16'hCD56, 16'hCD96, 16'hEE9B, 16'hF71D, 16'hF6DC, 16'hDE19, 16'hEE9B, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hE69A, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD618, 16'hA492, 16'h8BCF, 16'hDE59, 16'hDE59, 16'hAD13, 16'hB596, 16'hF79E, 16'h83CF, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'h734D, 16'hF79D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h83CF, 16'hEE9B, 16'hEEDC, 16'hEEDC, 16'hF71D, 16'hB514, 16'hC618, 16'hCE59, 16'h7B4E, 16'hE61A, 16'hC515, 16'hEE5A, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hEE9B, 16'h8A09, 16'hD556, 16'hFF5E, 16'hDE19, 16'hBCD4, 16'h49C8, 16'h000, 16'h2904, 16'h30C3, 16'h4144, 16'h000, 16'h730C, 16'hC555, 16'hD5D7, 16'h734C, 16'h000, 16'h1205, 16'h3AC8, 16'h4B0A, 16'h5B8C, 16'h5B8C, 16'h5B8C, 16'h5B8C, 16'h5B8C, 16'h5B8C, 16'h530A, 16'h4288, 16'h080, 16'h9C51, 16'hF71C, 16'hEEDC, 16'hFF5E, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hFF9F, 16'hEEDC, 16'hDE19, 16'hDDD8, 16'hCD96, 16'hCD96, 16'hCD96, 16'h4A07, 16'h2A06, 16'h5B8C, 16'h640E, 16'h640E, 16'h640E, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCC, 16'h5BCC, 16'h4B0A, 16'h0C1, 16'h1882, 16'h3903, 16'h4985, 16'h4986, 16'h2882, 16'h4144, 16'hEE9B, 16'hFF1E, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hE65A, 16'hEE5A, 16'hEE5A, 16'hEE5B, 16'hEE9B, 16'hF6DC, 16'hF6DD, 16'hEE9B, 16'h6A8A, 16'hAC10, 16'hCCD4, 16'hD556, 16'hCD96, 16'hE65A, 16'hF71D, 16'hF6DC, 16'hDE19, 16'hE65A, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hE69B, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hD5D8, 16'hACD3, 16'h628A, 16'hD618, 16'hDE59, 16'hBD55, 16'h9492, 16'hFFDF,
        16'h83CF, 16'hDE5A, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'h7B4E, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDF1B, 16'h8BD0, 16'hF6DC, 16'hEEDB, 16'hEEDB, 16'hF71D, 16'h9411, 16'hDEDB, 16'hCE59, 16'h7B4E, 16'hE619, 16'hCD56, 16'hEE5B, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D,
        16'hF71D, 16'hF71D, 16'hF6DC, 16'hA34E, 16'hE556, 16'hD5D7, 16'hC515, 16'h624A, 16'h000, 16'h3104, 16'h3103, 16'h2082, 16'h000, 16'h9C51, 16'hD5D7, 16'hD597, 16'h62CA, 16'h000, 16'h3287, 16'h4B0A, 16'h5B8C, 16'h63CD, 16'h63CD, 16'h5BCD, 16'h63CD, 16'h63CD, 16'h63CD, 16'h63CE, 16'h63CE, 16'h63CD, 16'h530B, 16'h000, 16'hA4D2, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hF71D, 16'hEE9B, 16'hACD3, 16'h000, 16'h4B0A, 16'h640D, 16'h640D, 16'h640E, 16'h640D, 16'h640E, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5B8C, 16'h5BCD, 16'h4B0B, 16'h040, 16'h4A07, 16'h4145, 16'h3842,
        16'h38C3, 16'h5186, 16'hEE9B, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hE65A, 16'hEE5A, 16'hEE5A, 16'hEE5B, 16'hEE9B, 16'hF6DC, 16'hFF1D, 16'hEE9B, 16'h6A8A, 16'hABD0, 16'hC4D4, 16'hCD56, 16'hCD56, 16'hDE19, 16'hF6DC, 16'hF6DC, 16'hDE19, 16'hE65A, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hE69B, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hBD55, 16'h3904, 16'hBD55, 16'hE659, 16'hCDD7, 16'h83D0, 16'hFFDF, 16'h9451, 16'hD619, 16'hEEDB, 16'hE69B, 16'hEEDC, 16'h8BD0, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h9C52, 16'hF71D, 16'hEEDB, 16'hEEDC, 16'hF6DC, 16'h838E, 16'hEF5D, 16'hCE59, 16'h834E, 16'hDDD8, 16'hD557, 16'hE65A, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hAC11, 16'hB3D0, 16'hC555, 16'h7B4D, 16'h000, 16'h2904, 16'h3904, 16'h30C3, 16'h000, 16'hAC92, 16'hD5D7, 16'hD5D7, 16'h8BCF, 16'h000, 16'h32C8, 16'h4B4B, 16'h63CD, 16'h5B8D, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h63CD, 16'h63CD, 16'h63CD, 16'h63CD, 16'h63CD, 16'h63CE, 16'h6C0E, 16'h634C, 16'h000, 16'hBD96, 16'hFFDF, 16'hFF5E, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF5F, 16'hFF5F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'h9452, 16'h0C0, 16'h5B8C, 16'h640E, 16'h63CD, 16'h63CE, 16'h5BCD, 16'h63CD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5B8D, 16'h5B8C, 16'h63CE, 16'h2246, 16'h5A89, 16'hC514, 16'h7ACB, 16'h3000, 16'h61C7, 16'hEE9B, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hE61A, 16'hEE5A, 16'hEE5A, 16'hEE5B, 16'hEE5B, 16'hF6DC, 16'hFF1D, 16'hEE9B, 16'h6249, 16'hAC10, 16'hC4D4, 16'hCD96, 16'hCD56, 16'hD5D8, 16'hF6DC, 16'hF6DC, 16'hDE19, 16'hE65A, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC,
        16'hEE9B, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hC596, 16'h3945, 16'h9C92, 16'hE659, 16'hD618, 16'h838E, 16'hFF9E, 16'hA514, 16'hCDD7, 16'hEEDC, 16'hE69B, 16'hEEDC, 16'hA492, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'hBD55, 16'hF71D, 16'hEE9B, 16'hF6DC, 16'hE69B, 16'h7B8E, 16'hFFDF, 16'hCE59, 16'h834E, 16'hDDD8, 16'hD597, 16'hE65A, 16'hEEDC, 16'hF6DD, 16'hF71D, 16'hF71D,
        16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1E, 16'hBCD4, 16'h9BCF, 16'h93D0, 16'h000, 16'h28C3, 16'h3903, 16'h3944, 16'h000, 16'hACD2, 16'hDE17, 16'hD5D7, 16'hBD55, 16'h2144, 16'h1A05, 16'h4B4A, 16'h63CD, 16'h5B8D, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h63CD, 16'h63CD, 16'h63CD, 16'h63CE, 16'h63CE, 16'h63CE, 16'h63CE, 16'h6C0E, 16'h530A, 16'h3185, 16'hEF1C, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hF75E, 16'h4A49, 16'h000, 16'h3B09, 16'h640D, 16'h640E, 16'h640E, 16'h63CD, 16'h640D, 16'h63CE, 16'h63CD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD,
        16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5B8C, 16'h6C0E, 16'h538B, 16'h080, 16'hBD14, 16'hDD97, 16'h9B8E, 16'h7248, 16'hF6DC, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hE61A, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hF6DC, 16'hFF1D, 16'hEE5A, 16'h6249, 16'hAC11, 16'hC4D4, 16'hD596, 16'hCD96, 16'hD597, 16'hF6DC, 16'hF6DC, 16'hDE5A, 16'hDE19, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hE69B, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hCDD7, 16'hC596, 16'h5289, 16'h7B4D, 16'hDE59, 16'hDE59, 16'h83CF, 16'hF75D, 16'hBD96, 16'hBD55, 16'hEEDC, 16'hE69B, 16'hEEDC, 16'hB515, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h8C10, 16'hD618, 16'hF6DC, 16'hEE9B, 16'hF6DC, 16'hD5D8, 16'h8C51, 16'hFFDF, 16'hD69A, 16'h838E, 16'hDDD8, 16'hD597, 16'hE65A, 16'hEEDC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1E, 16'hD5D8, 16'h6A8A, 16'h000, 16'h1841, 16'h30C3, 16'h4945, 16'h000, 16'h9C50, 16'hD617, 16'hCD96, 16'hD5D7, 16'h9C51, 16'h000, 16'h42C9, 16'h5B8D, 16'h5B8D, 16'h5BCD, 16'h63CD, 16'h63CD, 16'h63CD, 16'h63CD, 16'h5BCD, 16'h5BCD, 16'h63CD, 16'h63CD, 16'h63CD, 16'h63CE, 16'h63CE, 16'h63CE,
        16'h6C0E, 16'h182, 16'hB555, 16'hFFDF, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hF71D, 16'hAD14, 16'hAD55, 16'h9D14, 16'h640E, 16'h640E, 16'h640E, 16'h640E, 16'h640E, 16'h640E, 16'h5BCD, 16'h640E, 16'h6C0F, 16'h6C4F, 16'h644F, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h63CE, 16'h6C4F, 16'h5BCD, 16'h100, 16'h9C10, 16'hDD97, 16'h828A, 16'h82CB, 16'hF6DC, 16'hFF1D, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hE619, 16'hEE5A, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hF6DC, 16'hFF1D, 16'hE65A, 16'h6209, 16'hAC11,
        16'hC514, 16'hCD96, 16'hCD96, 16'hCD97, 16'hEE9B, 16'hF6DC, 16'hE65A, 16'hDE19, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hE69B, 16'hCE18, 16'hCE17, 16'hCE17, 16'hCDD7, 16'hC5D7, 16'h6B4C, 16'h5289, 16'hCDD7, 16'hDE5A, 16'h83CF, 16'hEF1C, 16'hCE59, 16'hACD4, 16'hEEDC, 16'hE69B, 16'hEEDC, 16'hC596, 16'h9451, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h7B8E, 16'hE65A, 16'hEEDC, 16'hEE9B, 16'hF71D,
        16'hBD56, 16'hAD14, 16'hFFDF, 16'hD65A, 16'h8B8F, 16'hCD56, 16'hD597, 16'hE65A, 16'hEE9B, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hFF1D, 16'hE65A, 16'h2881, 16'h000, 16'h3103, 16'h4945, 16'h800, 16'h7B0C, 16'hD5D7, 16'hCDD7, 16'hCD96, 16'hD5D7, 16'h83CE, 16'h140, 16'h538C, 16'h63CD, 16'h5BCD, 16'h5BCD, 16'h63CD, 16'h63CD, 16'h5BCD, 16'h63CD, 16'h63CD, 16'h63CD, 16'h63CD, 16'h63CD, 16'h63CD, 16'h640E, 16'h640E, 16'h63CE, 16'h63CE, 16'h4B0A, 16'h630B, 16'hF75E, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFFDF, 16'hFF9F,
        16'hFF9F, 16'h8CD2, 16'h5BCD, 16'h6C0E, 16'h640E, 16'h640E, 16'h640E, 16'h640E, 16'h6C4F, 16'h640E, 16'h640E, 16'h640F, 16'h644F, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h640E, 16'h640E, 16'h640E, 16'h6C4F, 16'h640D, 16'h1C0, 16'h8BCF, 16'hD556, 16'h4000, 16'h8B4D, 16'hFEDD, 16'hF71D, 16'hFF1D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hE619, 16'hEE5A, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hF6DC, 16'hFF1D, 16'hE65A, 16'h5A08, 16'hAC51, 16'hC515, 16'hCD96, 16'hCD96, 16'hCD56, 16'hE65A, 16'hF6DC, 16'hE65A, 16'hDE19, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hE69B, 16'hCE18, 16'hCE17, 16'hCE17, 16'hCDD7, 16'hC5D7, 16'h738C, 16'h3A06, 16'hBD55, 16'hE65A, 16'h83CF, 16'hDEDB, 16'hDEDB, 16'hA492, 16'hEEDC, 16'hE69B, 16'hEEDB, 16'hCDD7, 16'h8410, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h7B4E, 16'hEEDC, 16'hEEDC, 16'hEE9B, 16'hF71D, 16'hA493, 16'hC5D7, 16'hFFDF, 16'hD65A, 16'h8B8F, 16'hC515, 16'hCD56, 16'hEE5A, 16'hEE9B, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF6DD, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF71D, 16'hF6DC, 16'h7B4D, 16'h000, 16'h4185, 16'h30C2, 16'h4104, 16'hC555, 16'hD5D7, 16'hCD96, 16'hCD96, 16'hCDD7, 16'h630B, 16'h205, 16'h63CD, 16'h63CD, 16'h5BCD, 16'h5BCD,
        16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h63CD, 16'h63CD, 16'h63CD, 16'h63CD, 16'h63CD, 16'h63CE, 16'h63CE, 16'h63CD, 16'h63CE, 16'h6BCD, 16'h29C4, 16'hDE9A, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'h8CD2, 16'h5BCD, 16'h6C0E, 16'h640E, 16'h640E, 16'h640E, 16'h6C4F, 16'h6C4F, 16'h53CD, 16'h53CD, 16'h538D, 16'h5BCE, 16'h6C4F, 16'h640E, 16'h640E, 16'h640E, 16'h640E, 16'h640E, 16'h640F, 16'h640D, 16'h1C0, 16'h940F, 16'hC514, 16'h1800, 16'hA3CF, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D,
        16'hF71D, 16'hEE9C, 16'hDE19, 16'hEE5A, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hF6DC, 16'hFF1D, 16'hDE19, 16'h5187, 16'hAC51, 16'hC555, 16'hCD96, 16'hCD96, 16'hCD56, 16'hDE19, 16'hF6DC, 16'hE65A, 16'hDE19, 16'hEEDC, 16'hEEDC, 16'hEE9B, 16'hEEDC, 16'hEE9B, 16'hCE18, 16'hCE17, 16'hCE17, 16'hCE17, 16'hC5D7, 16'h7B8D, 16'h4A88, 16'h9C92, 16'hE69A, 16'h9410, 16'hD69A, 16'hEF1C, 16'h9C51, 16'hEEDC, 16'hE69B, 16'hEEDB, 16'hD618, 16'h7B8F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8C10, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'h9410, 16'hD659, 16'hFFDF, 16'hCE59, 16'h8B8F, 16'hBCD4, 16'hCD56, 16'hEE5A, 16'hEE5B, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hA451, 16'h000, 16'h2841, 16'h2800, 16'h9C0F, 16'hD5D7, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'h4A49, 16'h2A87, 16'h6C0E, 16'h63CD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h63CD, 16'h640E, 16'h6C0E, 16'h640E, 16'h6C0E, 16'h640E, 16'h63CD, 16'h63CE, 16'h6C0F, 16'h744F, 16'h740F, 16'h3246, 16'hB555, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hB556, 16'hB595, 16'hAD96, 16'h7C90, 16'h6C4F, 16'h6C0F, 16'h640E, 16'h640E, 16'h640F, 16'h640E, 16'h5C0E, 16'h4B8C, 16'h53CD, 16'h4B8C, 16'h434C, 16'h640F, 16'h6C4F, 16'h640E, 16'h640E, 16'h640E, 16'h640E, 16'h6C0E, 16'h63CD, 16'h201, 16'h9C50, 16'hAC51, 16'h000, 16'hAC51, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hEE9B, 16'hDDD9, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEEDC, 16'hFF1D, 16'hD5D8, 16'h4986, 16'hAC92, 16'hC555, 16'hCD96, 16'hCD96, 16'hC596, 16'hD618, 16'hF6DC, 16'hE65A, 16'hD619, 16'hEE9B, 16'hEEDC, 16'hEEDB, 16'hEEDC, 16'hEE9B, 16'hCE18, 16'hCE17, 16'hCE17, 16'hCDD7, 16'hCE17, 16'h7BCE, 16'h530A, 16'h83CF, 16'hE69A, 16'h9C52, 16'hCE59, 16'hEF5D, 16'h9410, 16'hEEDB, 16'hE69B, 16'hEEDB, 16'hDE19, 16'h7B8E, 16'hFF9F,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'hACD3, 16'hF6DC, 16'hEE9B, 16'hEEDC, 16'hEEDC, 16'h838E, 16'hE6DB, 16'hFFDF, 16'hCE59, 16'h8B8F, 16'hBCD3, 16'hCD56, 16'hEE5A, 16'hE65A, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1E, 16'hC555, 16'h000, 16'hA451, 16'h834D,
        16'hA451, 16'hD5D7, 16'hCD96, 16'hCD96, 16'hCD96, 16'hC596, 16'h4A48, 16'h2287, 16'h6C0E, 16'h63CD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h640E, 16'h640E, 16'h63CE, 16'h5BCD, 16'h6C0E, 16'h6C0F, 16'h6C0E, 16'h744F, 16'h7450, 16'h7450, 16'h7C50, 16'h4B0A, 16'h9C51, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'h7B8E, 16'h204, 16'h7490, 16'h8D53, 16'h8D53, 16'h8512, 16'h84D2, 16'h7490, 16'h640E, 16'h6450, 16'h6C50, 16'h644F, 16'h644F, 16'h5C0F, 16'h6450, 16'h6C90, 16'h6C4F, 16'h640E, 16'h640E, 16'h640E, 16'h640E, 16'h6C0E, 16'h63CD, 16'h244, 16'h940F, 16'h82CB, 16'h3800, 16'hBCD4, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D,
        16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hEE9B, 16'hDDD8, 16'hEE9B, 16'hE65B, 16'hEE5B, 16'hEE5A, 16'hEEDC, 16'hFF1D, 16'hCD97, 16'h4986, 16'hAC92, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hD5D8, 16'hEEDC, 16'hE69A, 16'hD5D8, 16'hEE9B, 16'hEE9B, 16'hEEDB, 16'hEEDC, 16'hE69B, 16'hCE18, 16'hC657, 16'hCE17, 16'hC617, 16'hCE17, 16'h7BCE, 16'h638C, 16'h62CB, 16'hDE19, 16'hACD4, 16'hC5D7, 16'hF79E, 16'h8BD0, 16'hEEDB, 16'hE69B, 16'hEEDB, 16'hDE59, 16'h7B8E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'hBD56, 16'hF6DC, 16'hEE9B, 16'hEEDC, 16'hE65A, 16'h7B8E, 16'hEF5D, 16'hFFDF, 16'hD65A, 16'h8B8F, 16'hB493, 16'hCD56, 16'hEE5B, 16'hE65A, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF6DC, 16'hEE9C, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hFF1D, 16'hD5D8, 16'h8B4D, 16'hD596, 16'h40C3, 16'hA451, 16'hD5D7, 16'hCD96, 16'hCD96, 16'hCD96, 16'hBD55, 16'h3A06, 16'h2AC7, 16'h538C, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h640E, 16'h640E, 16'h63CD, 16'h5BCD, 16'h538C, 16'h5BCD, 16'h63CE, 16'h6C4F, 16'h744F, 16'h744F, 16'h7C90, 16'h7C90, 16'h63CD, 16'h7B8E, 16'hFF5E, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hA4D3, 16'h3288, 16'h84D2, 16'h8D53, 16'h8D13, 16'h8513, 16'h8513, 16'h7CD2, 16'h7CD2, 16'h8D95, 16'h8D95, 16'h8D95, 16'h8D95, 16'h8D94, 16'h8553, 16'h8554, 16'h74D1, 16'h640E, 16'h640D, 16'h63CE, 16'h640E, 16'h6C0E, 16'h5BCC, 16'h2286, 16'h9C0F, 16'h7249, 16'hA34D, 16'hCD56, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hF71D, 16'hEE5B, 16'hDDD8, 16'hEE9B, 16'hEE5B, 16'hE65B, 16'hEE5B, 16'hF6DC, 16'hFF1D, 16'hC556, 16'h4985, 16'hAC92, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCDD7, 16'hEEDC, 16'hE69A, 16'hD5D8, 16'hEE9B, 16'hEE9B, 16'hEEDB, 16'hEEDC, 16'hE69B, 16'hCE18, 16'hC657, 16'hC617, 16'hC617, 16'hCE18, 16'h7BCE, 16'h6B8C,
        16'h528A, 16'hD619, 16'hB515, 16'hB596, 16'hF79E, 16'h83CF, 16'hE69B, 16'hE69B, 16'hEEDB, 16'hDE5A, 16'h7B8E, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h8C11, 16'hCDD8, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hDE59, 16'h83CF, 16'hF79E, 16'hFFDF, 16'hD69A, 16'h93D0, 16'hAC52, 16'hC556, 16'hEE5B, 16'hDE19, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF71D, 16'hF71D,
        16'hF71D, 16'hFF1D, 16'hF6DD, 16'hEE9B, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF71D, 16'hEE9B, 16'h938E, 16'hAC51, 16'h000, 16'h938E, 16'hD5D7, 16'hCD96, 16'hC555, 16'hC555, 16'hD619, 16'hE6DB, 16'hEF5D, 16'hCE59, 16'h534C, 16'h63CE, 16'h5BCD, 16'h5BCD, 16'h5BCD, 16'h640E, 16'h5C0D, 16'h5BCD, 16'h5BCD, 16'h538C, 16'h63CE, 16'h6C0E, 16'h744F, 16'h7C90, 16'h744F, 16'h744F, 16'h7C90, 16'h744F, 16'h6B0B, 16'hF71D, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hBD96, 16'h1206, 16'h8512, 16'h8D53, 16'h8D53, 16'h8512, 16'h8513, 16'hA617, 16'hAE58, 16'h9595, 16'h9595, 16'h9595, 16'h8D95, 16'h9595, 16'h9595, 16'h7D13, 16'h6450, 16'h5C0E, 16'h7491, 16'h7490, 16'h6C0F, 16'h640E,
        16'h4B8B, 16'h4AC9, 16'h938E, 16'hA38F, 16'hC452, 16'hCD97, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hEE5A, 16'hDDD8, 16'hEE9B, 16'hEE5B, 16'hE65B, 16'hEE5B, 16'hF6DC, 16'hFF1D, 16'hBD15, 16'h51C7, 16'hAC93, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hEE9B, 16'hE69B, 16'hD5D8, 16'hEE9B, 16'hEE9B, 16'hEEDB, 16'hEEDC, 16'hE69B, 16'hCE58, 16'hCE17, 16'hCE17, 16'hC617, 16'hCE18, 16'h83CF, 16'h638C, 16'h5ACB, 16'hD619, 16'hBD56, 16'hB555, 16'hF79E, 16'h83CF, 16'hE6DB, 16'hE69B, 16'hEEDB, 16'hDE59, 16'h7B8E, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h83CF, 16'hE65A, 16'hEEDC, 16'hEEDB, 16'hEE9B, 16'hD619, 16'h8C51, 16'hFFDF, 16'hFFDF, 16'hD69B, 16'h9BD0, 16'hAC52, 16'hCD56, 16'hEE9B, 16'hDE19, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hEE5B, 16'hF6DC, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'h9C10, 16'h6A48, 16'h3800, 16'h7249, 16'hCD55, 16'hC555, 16'hD618, 16'hEF1C, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hF79D, 16'h5BCD, 16'h53CD, 16'h538D, 16'h53CD, 16'h5BCD, 16'h6C4F, 16'h640E, 16'h640E, 16'h6C4F, 16'h7490, 16'h8512, 16'h8D12, 16'h8D13, 16'h8D53, 16'h7C91, 16'h8C91, 16'h8CD2, 16'h8490, 16'h630A, 16'hEEDC, 16'hFF9F, 16'hFF5E, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hD65A, 16'h19C5, 16'h84D2, 16'h8D54, 16'h8512, 16'h9554, 16'hB658, 16'hBE99, 16'hB699, 16'hAE17, 16'h8D54, 16'h9595, 16'h9595, 16'h9595, 16'h8D94, 16'h9594, 16'hDF1C, 16'hD71B, 16'h7CD1, 16'h7CD2, 16'h8513, 16'h84D2, 16'h3B4A, 16'h83CE, 16'h938E, 16'hCCD4, 16'hBC11, 16'hDE18, 16'hFF5E, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hE61A, 16'hDDD9, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hFF1D, 16'hAC93, 16'h5207, 16'hB4D3, 16'hCD97, 16'hCD96, 16'hCD96, 16'hCD96, 16'hCD96, 16'hE69A, 16'hE69B, 16'hCDD8,
        16'hE69B, 16'hEEDB, 16'hEEDB, 16'hEEDB, 16'hE69B, 16'hCE58, 16'hC618, 16'hC618, 16'hC617, 16'hCE58, 16'h840F, 16'h638C, 16'h5ACA, 16'hD5D9, 16'hC556, 16'hAD55, 16'hF79E, 16'h83CF, 16'hE69B, 16'hE69B, 16'hEEDB, 16'hDE59, 16'h7BCF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h83CF, 16'hEEDC, 16'hEEDC, 16'hEE9B, 16'hE69B, 16'hD5D8, 16'h9492, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h9C10, 16'hB492, 16'hCD56, 16'hEE9B,
        16'hDE19, 16'hE65B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hEE5B, 16'hF69C, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hFF1E, 16'hBD14, 16'h2000, 16'h4083, 16'h4840, 16'hBCD3, 16'hEEDB, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hD699, 16'h8D12, 16'h53CD, 16'h6450, 16'h74D1, 16'h7D12, 16'h7D12, 16'h8513, 16'h7450, 16'h7450, 16'h8D13, 16'h8D13, 16'h8D53, 16'h8D13, 16'h9554, 16'h8D13, 16'hBE59, 16'hF79E, 16'hCE59, 16'h94D2, 16'h6B0B, 16'hEEDC, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hF71D, 16'h5B0B, 16'h7C91, 16'h8D53, 16'h8D54, 16'hB699, 16'hBE99, 16'hB699, 16'hB699, 16'hB699,
        16'hA617, 16'h8D54, 16'h8D54, 16'h9595, 16'h9DD6, 16'hB659, 16'hD6DB, 16'hDF1C, 16'hAE18, 16'h8D54, 16'h8513, 16'h8D53, 16'h2B09, 16'hACD2, 16'h9B8E, 16'hE557, 16'hABCF, 16'hEE9A, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hE619, 16'hDE19, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hFF1D, 16'hA452, 16'h6289, 16'hB4D4, 16'hCD97, 16'hCD96, 16'hCD96, 16'hCD96, 16'hC596, 16'hE65A, 16'hE69B, 16'hCDD8, 16'hE69B, 16'hEEDB, 16'hEE9B, 16'hEEDB, 16'hE69B, 16'hC658, 16'hC658, 16'hC658, 16'hC617, 16'hCE58, 16'h840F, 16'h5B4B, 16'h5289, 16'hD619, 16'hC556, 16'hA514, 16'hF79E, 16'h83CF, 16'hEEDB, 16'hE69B, 16'hEEDB, 16'hD619, 16'h83CF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9B, 16'h83CF, 16'hF6DC, 16'hEEDC, 16'hE69B, 16'hE69B, 16'hC597, 16'hA4D3, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h9C11, 16'hB492, 16'hCD56, 16'hEE9B, 16'hDE19, 16'hE65A, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hFF1D, 16'hF69C, 16'hEE5B, 16'hFF1D, 16'hF6DD, 16'hF6DD, 16'hFF1E, 16'hD5D8, 16'h48C0, 16'h8B0C, 16'h2000, 16'hBD14, 16'hFFDF, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'h5B0B, 16'h246, 16'h7D12, 16'h8D94, 16'h8D94, 16'h8D54, 16'h8554, 16'h8513, 16'h8513, 16'h8D13, 16'h8513, 16'h8D54, 16'h8D54,
        16'h9554, 16'h9554, 16'h9D95, 16'hBE58, 16'hBE99, 16'hBE58, 16'hB616, 16'h734C, 16'hE69B, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hA4D3, 16'h5BCD, 16'h9D95, 16'hB699, 16'hB699, 16'hB699, 16'hB699, 16'hB699, 16'hB659, 16'hBE9A, 16'hBE9A, 16'hB659, 16'hAE18, 16'hB659, 16'hB699, 16'hB659, 16'hAE59, 16'hBE9A, 16'hB659, 16'h8D14, 16'h7CD1, 16'h73CD, 16'hC555, 16'hBC52, 16'hED97, 16'hA38F, 16'hFEDC, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hE619, 16'hE619, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hF6DC,
        16'hF6DC, 16'h8B8F, 16'h6ACB, 16'hB514, 16'hCDD7, 16'hCD96, 16'hCD96, 16'hCD96, 16'hC596, 16'hDE59, 16'hE69B, 16'hCDD8, 16'hE69A, 16'hEEDB, 16'hE69B, 16'hEE9B, 16'hE69A, 16'hCE58, 16'hC658, 16'hC658, 16'hC657, 16'hCE58, 16'h8C50, 16'h5B0A, 16'h62CB, 16'hDE1A, 16'hBD56, 16'hA514, 16'hEF5D, 16'h838F, 16'hE6DB, 16'hE69B, 16'hEEDB, 16'hCE18, 16'h8C10, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h9451, 16'hF71D,
        16'hEEDB, 16'hE69B, 16'hEE9B, 16'hC596, 16'hB555, 16'hFFDF, 16'hFFDF, 16'hDEDA, 16'hA451, 16'hAC51, 16'hCD97, 16'hEE9B, 16'hE65A, 16'hDE19, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF6DC, 16'hDE19, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF6DC, 16'h6A89, 16'hD4D4, 16'hABD0, 16'h5943, 16'hF71C, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hFF9F, 16'hA4D3, 16'h1C4, 16'h74D1, 16'h8D94, 16'h8554, 16'h8554, 16'h8553, 16'h8513, 16'hA617, 16'hB659, 16'h9DD6, 16'h8D54, 16'h8D54, 16'h8D54, 16'h9554, 16'hAE57, 16'hB658, 16'hB658, 16'hB658, 16'hBE58, 16'h83CE, 16'hE6DC, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E,
        16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hDE9B, 16'h534B, 16'h9595, 16'hBE99, 16'hB699, 16'hB69A, 16'hB699, 16'hB699, 16'hC6DB, 16'hD71D, 16'hDF5E, 16'hDF5E, 16'hD71D, 16'hC69A, 16'hB659, 16'hBE99, 16'hBE9A, 16'hB69A, 16'hB65A, 16'hA5D7, 16'h4BCC, 16'hBD55, 16'hC4D4, 16'hE556, 16'hDD15, 16'hB452, 16'hFF1D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF71D, 16'hEEDC, 16'hF6DC, 16'hF6DD, 16'hF71D, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hDDD9, 16'hE619, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hF6DC, 16'hEE9B, 16'h6ACB, 16'h730C, 16'hBD14, 16'hCDD7, 16'hCD96, 16'hCD96, 16'hCD96, 16'hC596, 16'hDE19, 16'hE69B, 16'hCDD8, 16'hDE5A, 16'hEEDB, 16'hE69B, 16'hEE9B, 16'hE69A, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hCE58, 16'h8C50, 16'h4247, 16'h7B8E, 16'hE65A, 16'hBD56, 16'hAD55, 16'hEF5D, 16'h83CF, 16'hEEDB, 16'hE69B, 16'hEEDC, 16'hC596, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC5D7, 16'hA492, 16'hF71D, 16'hEE9B, 16'hE69A, 16'hEEDB, 16'hBD55, 16'hB556, 16'hFFDF, 16'hFFDF, 16'hDEDA, 16'hAC52, 16'hA411, 16'hCD96, 16'hEE9B, 16'hE65A, 16'hD5D8, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hFF1D, 16'hE619, 16'hEE9B, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hFF1D, 16'h9C10, 16'hA34E, 16'hF5D8, 16'h930C, 16'hAC92, 16'hFFDF, 16'hFF9E, 16'hFF5E, 16'hFF9F, 16'hDE5A,
        16'h182, 16'h644F, 16'h8554, 16'h8D94, 16'h8554, 16'h8D54, 16'hA618, 16'hB699, 16'hB659, 16'hB69A, 16'hAE58, 16'hAE18, 16'hBE59, 16'hBE99, 16'hAE17, 16'hAE17, 16'hB658, 16'hB658, 16'hBE58, 16'h8C50, 16'hEF1D, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFFDF, 16'hA555, 16'h6C50, 16'hAE58, 16'hB69A, 16'hB699, 16'hBE9A, 16'hD71D, 16'hDF5E, 16'hD71E, 16'hCEDC, 16'hCF1C, 16'hDF5E, 16'hDF1E, 16'hCEDC, 16'hBE9A, 16'hB65A, 16'hB65A, 16'hBE9B, 16'h9DD6, 16'h8450, 16'hE65A, 16'hCC93, 16'hFDD9, 16'hBC11, 16'hC555, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF6DD, 16'hF6DC, 16'hEE9C, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF6DD, 16'hF6DC, 16'hF6DC,
        16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hDDD8, 16'hE61A, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hF6DC, 16'hE65A, 16'h5208, 16'h834D, 16'hC555, 16'hCDD7, 16'hCD96, 16'hCD96, 16'hCD96, 16'hC596, 16'hD618, 16'hE69B, 16'hCDD8, 16'hDE5A, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hE69A, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hCE58, 16'h8C51, 16'h1982, 16'h8C10, 16'hE69B, 16'hB515, 16'hB596, 16'hE71C, 16'h83CF, 16'hEEDB, 16'hE69A, 16'hEEDC, 16'hACD3, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB555, 16'hAD14, 16'hF71C, 16'hE69B, 16'hE69A, 16'hEEDC, 16'hB555, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'hAC92, 16'hAC51, 16'hCD97, 16'hEE9B, 16'hE65A, 16'hD5D8, 16'hEE9B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hFF1D, 16'hEE5B, 16'hE619, 16'hFF1D, 16'hF6DD, 16'hF6DD, 16'hFF1D, 16'hD5D8, 16'h6945, 16'hDD15, 16'hF65A, 16'hAC11, 16'hD5D8, 16'hFF9F, 16'hFF5E, 16'hFF9E, 16'hFF9F, 16'h7BCF, 16'h330A, 16'h8554, 16'h8554, 16'h8D94, 16'hAE58, 16'hB699, 16'hB699, 16'hB699, 16'hB659, 16'hCEDC, 16'hDF5E, 16'hDF5E, 16'hDF5E, 16'hD71C, 16'hBE99, 16'hB658, 16'hAE18, 16'hB658, 16'hB555, 16'hFF5E, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFFDF, 16'hF79E, 16'h8C92, 16'h9555, 16'hBEDB, 16'hC6DC, 16'hD71D, 16'hDF5E, 16'hDF5E, 16'hDF1E, 16'hB65A, 16'hBE9B, 16'hDF5E, 16'hDF1D, 16'hDF5E, 16'hD71D, 16'hBE9A, 16'hBE9A, 16'hBE9A, 16'h7450, 16'hE6DB, 16'hF69B, 16'hE556, 16'hF5D8, 16'hBBD0, 16'hE619, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hEE9C, 16'hEEDC, 16'hF6DD, 16'hF6DD, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hD597, 16'hE65A, 16'hEE5B, 16'hE65B, 16'hE65B, 16'hE65A, 16'hF6DC, 16'hDE19, 16'h4185, 16'h8BCF, 16'hC596, 16'hCDD7, 16'hCD96, 16'hCD96, 16'hCD96, 16'hC596, 16'hD5D7, 16'hE69A, 16'hCE18, 16'hDE59, 16'hEE9B, 16'hE69B, 16'hEE9B, 16'hDE9A, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hCE58, 16'h8C51, 16'h000, 16'hACD3, 16'hEE9B, 16'hB514, 16'hB596, 16'hE71C, 16'h8C10, 16'hEEDC, 16'hE69A,
        16'hEEDC, 16'h9411, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA4D3, 16'hBD55, 16'hF71C, 16'hE69B, 16'hE69B, 16'hEEDC, 16'hB515, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'hAC92, 16'hA451, 16'hCD96, 16'hEE9B, 16'hEE5B, 16'hD5D8, 16'hE65B, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hF6DC, 16'hDDD8, 16'hF6DC, 16'hF6DD,
        16'hF6DD, 16'hF6DD, 16'hFEDD, 16'h830C, 16'hB3D0, 16'hEE19, 16'hFEDD, 16'hB493, 16'hF6DC, 16'hFF9F, 16'hFF5E, 16'hFFDF, 16'hD659, 16'h140, 16'h7D12, 16'h8D95, 16'hAE59, 16'hB699, 16'hB659, 16'hB699, 16'hB699, 16'hBE9A, 16'hD75E, 16'hDF5E, 16'hCF1C, 16'hC6DC, 16'hDF5E, 16'hDF5E, 16'hD71D, 16'hCEDC, 16'hBE59, 16'hD659, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFFDF, 16'hDEDB, 16'h9D96, 16'hC71C, 16'hD75E, 16'hDF5E, 16'hDF5E, 16'hDF5E, 16'hDF5E, 16'hC6DC, 16'hC6DC, 16'hDF1E, 16'hDF1D, 16'hDF1D, 16'hDF5E, 16'hD71C, 16'hC6DB, 16'h7CD2, 16'hCE59, 16'hFF9F, 16'hEDD8, 16'hF597, 16'hED57, 16'hABCF, 16'hF69C, 16'hF71D, 16'hF6DD, 16'hF6DD,
        16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hE65B, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hEEDC, 16'hEE9C, 16'hF6DC, 16'hEE9B, 16'hD597, 16'hEE5A, 16'hE69B, 16'hE65B, 16'hE65B, 16'hE65A, 16'hF6DC, 16'hCD97, 16'h000, 16'h9410, 16'hCD97, 16'hCD97, 16'hCD97, 16'hCD96, 16'hCD96, 16'hC596, 16'hCDD7, 16'hE69A, 16'hCE18, 16'hD659, 16'hE69B, 16'hE69B, 16'hE69B, 16'hDE9A, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'h8450, 16'h000, 16'hBD96, 16'hEEDC, 16'hACD4, 16'hBDD7, 16'hDEDB, 16'h9451, 16'hEEDC, 16'hE69B, 16'hE69B, 16'h734D, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h8C51, 16'hC5D7, 16'hEEDC, 16'hE69B, 16'hE69B, 16'hEEDC, 16'hB515, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'hA492, 16'hAC92, 16'hCD56, 16'hEE9C, 16'hEE9B, 16'hDE18, 16'hE619, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hDDD8, 16'hE65A, 16'hFF1D, 16'hF6DD, 16'hF6DD, 16'hFF1E, 16'hC515, 16'h8209, 16'hE556, 16'hFEDC, 16'hF6DC, 16'hDE19, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'h8410, 16'h3B4B, 16'h9E17, 16'hB69A, 16'hB699, 16'hB699, 16'hB699, 16'hBE9A, 16'hD71D, 16'hDF5D, 16'hDF1D, 16'hC6DD, 16'h9E1A, 16'hCF1D, 16'hDF5E, 16'hDF5E, 16'hDF5E, 16'hC69A, 16'hE6DC, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFFDF, 16'hD69A, 16'hB659, 16'hC6DB, 16'hD71D, 16'hE79F, 16'hEF9F, 16'hEF9F, 16'hEF9F, 16'hE79F, 16'hE75E, 16'hDF5E, 16'hDF5E, 16'hDF1E, 16'hD71D, 16'hBE9A, 16'hC659, 16'hFF9F, 16'hF69C, 16'hED57, 16'hF5D8, 16'hD4D4, 16'hA3D0, 16'hFF1D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hFF1D, 16'hEE9B, 16'hEE9B, 16'hF71D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hF6DC, 16'hEE5B, 16'hD597, 16'hEE5B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hE65A, 16'hF6DC, 16'hB4D4, 16'h20C0, 16'hA491, 16'hCDD7, 16'hCD96, 16'hCDD7, 16'hCD96, 16'hC596, 16'hC596, 16'hCDD7, 16'hE69A, 16'hCE18, 16'hD659, 16'hE69B, 16'hE69B, 16'hE69B, 16'hDE9A, 16'hC658, 16'hC658, 16'hC658,
        16'hC658, 16'hCE98, 16'h7C0F, 16'h1881, 16'hD659, 16'hEEDC, 16'hA492, 16'hC618, 16'hD69A, 16'hA4D3, 16'hEEDC, 16'hE69B, 16'hD659, 16'h7BCE, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h8410, 16'hCDD8, 16'hEEDC, 16'hE69B, 16'hE69B, 16'hEEDC, 16'hAD14, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'hAC93, 16'hAC93, 16'hCD56, 16'hEE9B, 16'hEE9B, 16'hE619, 16'hDE19, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hEEDC, 16'hEEDC,
        16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hEE5A, 16'hD556, 16'hFEDD, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF69C, 16'h7A8B, 16'hB3CF, 16'hF65A, 16'hFF5E, 16'hF6DC, 16'hF71D, 16'hFF9F, 16'hFF9E, 16'hFF9F, 16'hEF1D, 16'h4B0A, 16'h5C4F, 16'hAE58, 16'hB699, 16'hB659, 16'hB69A, 16'hCF1C, 16'hDF5E, 16'hDF1D, 16'hDF1D, 16'hD71E, 16'hBEDC, 16'hD71E, 16'hE75E, 16'hDF5E, 16'hD71C, 16'hCE9A, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hDF1C, 16'hCEDB, 16'hCEDC, 16'hCF1C, 16'hD75D, 16'hDF5E, 16'hDF5E, 16'hE75E, 16'hE79F, 16'hE79F, 16'hD75E, 16'hD75E, 16'hC6DB,
        16'hB658, 16'hCE9A, 16'hEE9C, 16'hF65A, 16'hED57, 16'hFDD8, 16'hB3CF, 16'hBD15, 16'hFF1E, 16'hF6DD, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hE61A, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hE61A, 16'hD597, 16'hEE9B, 16'hE65A, 16'hEE5B, 16'hEE5B, 16'hE65A, 16'hF6DC, 16'hA452, 16'h3102, 16'hB513, 16'hCDD7, 16'hCD96, 16'hCDD7, 16'hCD96, 16'hC596, 16'hC596, 16'hCDD7, 16'hDE5A, 16'hCE18, 16'hD658, 16'hE69B, 16'hE69B, 16'hE69B, 16'hDE9A, 16'hC658, 16'hC698, 16'hC658, 16'hC658, 16'hCE99, 16'h73CE, 16'h5A8A, 16'hE69B, 16'hEEDB, 16'h9410, 16'hD6DA, 16'hCE58, 16'hB514, 16'hEEDB, 16'hEEDC, 16'hBD56, 16'h9492, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h738E, 16'hD618, 16'hEEDC, 16'hE69B, 16'hE69B, 16'hEEDC, 16'hACD4, 16'hC617, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hAC93, 16'hA492, 16'hC556, 16'hEE9B, 16'hEE5B, 16'hE65A, 16'hDDD8, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hD516, 16'hD597, 16'hFF1E, 16'hF71D, 16'hF71D, 16'hFF1E, 16'hC515, 16'h6800, 16'hDD57, 16'hFF1E, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF9F, 16'hFF9E, 16'hFFDF, 16'hEF1C, 16'h744F, 16'h7512, 16'hB69A, 16'hBE9A, 16'hCF1C, 16'hDF5E, 16'hDF5D, 16'hDF5D, 16'hDF5D, 16'hE75E, 16'hE79E, 16'hF7DF, 16'hEFDF, 16'hD71D, 16'hCE9A, 16'hEF5C, 16'hFF9F,
        16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hF75E, 16'hEF1D, 16'hE71D, 16'hDF1D, 16'hD71D, 16'hEF9E, 16'hD71C, 16'hAE58, 16'hAE99, 16'h9E16, 16'hBED9, 16'hEFDF, 16'hDEDC, 16'hE69B, 16'hFEDD, 16'hF65A, 16'hF597, 16'hF598, 16'h9B4D, 16'hE619, 16'hFF1D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hFF1D, 16'hE61A, 16'hEE9B, 16'hF71D, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hEEDC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hE619, 16'hD598, 16'hEE9B, 16'hE65A, 16'hEE5B, 16'hE65A, 16'hE65A, 16'hF69C, 16'h838F, 16'h49C6, 16'hB554, 16'hCDD7, 16'hCD96, 16'hC596, 16'hC596, 16'hC596,
        16'hC596, 16'hC597, 16'hDE59, 16'hCE58, 16'hCE18, 16'hE69A, 16'hE69B, 16'hE69B, 16'hD699, 16'hBE58, 16'hC698, 16'hC698, 16'hC658, 16'hCE98, 16'h634C, 16'h9451, 16'hEEDB, 16'hE69B, 16'h838F, 16'hE71C, 16'hB595, 16'hBD96, 16'hEEDB, 16'hEEDC, 16'h9411, 16'hC617, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h734D, 16'hDE59, 16'hEEDB, 16'hE69B, 16'hE69B, 16'hEEDC, 16'hACD4, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hE71C,
        16'hA492, 16'hAC93, 16'hC556, 16'hEE9C, 16'hE65B, 16'hE65A, 16'hD5D8, 16'hEE9B, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hEE19, 16'hA34E, 16'hCD97, 16'hFF5E, 16'hF71D, 16'hFF1D, 16'hF6DC, 16'h7A49, 16'hA34E, 16'hFEDD, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hF79E, 16'hDF1C, 16'h8513, 16'h8D95, 16'hC6DB, 16'hD75D, 16'hDF5E, 16'hE75E, 16'hE75E, 16'hE75E, 16'hE75E, 16'hEF9E, 16'hE75D, 16'hD71C, 16'hD6DB, 16'hEF1D, 16'hFF9F, 16'hFF9E, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1D,
        16'hFF1D, 16'hFF1D, 16'hFEDD, 16'hFF1D, 16'hDEDB, 16'hE75C, 16'hFFDF, 16'hE79D, 16'hE75D, 16'hE75C, 16'hBE58, 16'hC659, 16'hEE9B, 16'hFEDD, 16'hFEDD, 16'hF5D9, 16'hF5D8, 16'hDCD4, 16'h9B8F, 16'hFF1D, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DD, 16'hFF1D, 16'hEE9B, 16'hDDD8, 16'hF71D, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hDDD8, 16'hDDD8, 16'hEE9B, 16'hE65A, 16'hE65B, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'h6ACB, 16'h62CA, 16'hC595, 16'hCDD7, 16'hC596, 16'hC596, 16'hC596, 16'hC596, 16'hC596, 16'hC596, 16'hD659, 16'hCE58, 16'hCE18, 16'hDE9A, 16'hE69B, 16'hE69B, 16'hCE59, 16'hBE58, 16'hC698, 16'hC698, 16'hC698, 16'hC698, 16'h634C, 16'hBD96, 16'hEEDB, 16'hE69A, 16'h83CF, 16'hEF5D, 16'h9CD2, 16'hCDD7, 16'hEEDB, 16'hE69A, 16'h6B0C, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h734D, 16'hDE9A, 16'hEEDB, 16'hE69B, 16'hE69B, 16'hEEDC, 16'hACD4, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h9C92, 16'hACD3, 16'hC556, 16'hEE9C, 16'hE65B, 16'hEE9B, 16'hD5D8, 16'hE65A, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hEE9B, 16'hC494, 16'h5146, 16'hD5D8, 16'hFF5E, 16'hF6DD, 16'hFF5E, 16'hD597, 16'h4000, 16'hE5D8, 16'hFF1D, 16'hFEDC, 16'hFEDC, 16'hFF1D, 16'hFF9E, 16'hEF5D, 16'hBE59, 16'hB659, 16'hBF1B, 16'hAE59, 16'h9617, 16'hA659,
        16'hCF1C, 16'hDF5D, 16'hDF5D, 16'hD71C, 16'hD71C, 16'hD6DB, 16'hDF1C, 16'hEF5D, 16'hF75E, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5F, 16'hFF5F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1D, 16'hFEDD, 16'hFEDD, 16'hFF1D, 16'hEE5A, 16'hA515, 16'hE79E, 16'hDF5D, 16'hDEDB, 16'hDE5A, 16'hF6DC, 16'hEE5A, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hF5D8, 16'hFDD8, 16'hAB8E, 16'hC515, 16'hFF1E, 16'hF6DD, 16'hF71D, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hCD15, 16'hF69C, 16'hF6DD, 16'hF6DC, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF69C, 16'hD557, 16'hDE19, 16'hEE9B, 16'hE65A,
        16'hE65B, 16'hE65A, 16'hEE9B, 16'hE659, 16'h4186, 16'h838E, 16'hC5D6, 16'hC5D6, 16'hC596, 16'hC596, 16'hC596, 16'hC596, 16'hC596, 16'hC596, 16'hD618, 16'hCE58, 16'hCE18, 16'hDE5A, 16'hE69B, 16'hE69B, 16'hCE59, 16'hBE58, 16'hC698, 16'hC698, 16'hC698, 16'hBE57, 16'h528A, 16'hD618, 16'hEEDB, 16'hDE59, 16'h8C51, 16'hF79E, 16'h8410, 16'hCE18, 16'hEEDC, 16'hBD55, 16'h8C51, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hF79E, 16'h734D, 16'hDE9A, 16'hEEDB, 16'hE69B, 16'hE69B, 16'hEEDC, 16'hAD14, 16'hC617, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h9451, 16'hAD14, 16'hBD15, 16'hF69C, 16'hE65B, 16'hEE9B, 16'hDE19, 16'hDE19, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hD556, 16'h6208, 16'h20C1, 16'hD618, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'h8B4E, 16'hA38F, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hFEDD, 16'hF69B, 16'hBD96, 16'hEFDE, 16'hDF9E, 16'hC71C, 16'hCF5D, 16'hC71C, 16'hCF5D, 16'hCF9D, 16'hC75C, 16'hC71C, 16'hBE59, 16'hEF5D, 16'hF75E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hEE9B, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hFEDD, 16'hFEDD, 16'hFEDC, 16'hFEDD, 16'hBD56, 16'h9E17, 16'hC6DA, 16'hD659, 16'hEE9B, 16'hFE9C, 16'hFE9C, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hF5D9, 16'hE556, 16'h8B0D, 16'hF69C, 16'hFF1D, 16'hF6DD, 16'hF6DD, 16'hFEDD, 16'hFEDD, 16'hBC94, 16'hDE18, 16'hFF1D, 16'hF6DC, 16'hF71D, 16'hF6DD, 16'hF6DC, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hD557, 16'hE65A, 16'hEE5B, 16'hE65A, 16'hE65B, 16'hE65A, 16'hEE9B, 16'hD597, 16'h000, 16'h9451, 16'hCDD7, 16'hC596, 16'hC5D6, 16'hC5D6, 16'hC596, 16'hC596, 16'hC5D6, 16'hC596, 16'hCE18, 16'hCE58, 16'hCE18, 16'hD659, 16'hE69B, 16'hE69A, 16'hC658, 16'hBE58, 16'hC698, 16'hC698, 16'hC699, 16'hB5D6, 16'h630B, 16'hDE9A, 16'hEEDB, 16'hBD96, 16'h9CD3, 16'hF79E, 16'h738D, 16'hDE5A, 16'hEEDB, 16'h734D, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h734D, 16'hE69A, 16'hE6DB, 16'hE69B, 16'hE69B, 16'hEEDC, 16'hAD14, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9451, 16'hAD13, 16'hB4D4, 16'hF69C, 16'hE65B, 16'hEE5B, 16'hE61A, 16'hDDD8, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hDD98, 16'h82CC, 16'h52CA, 16'h28C2, 16'hBD55, 16'hFF1D, 16'hFF5F, 16'hE65A, 16'h4000,
        16'hDDD8, 16'hFEDD, 16'hF6DC, 16'hFEDC, 16'hFE9C, 16'hCDD7, 16'hCF1B, 16'hC6DB, 16'hDF5D, 16'hD6DB, 16'hF75D, 16'hEF5D, 16'hE79E, 16'hEF9E, 16'hEF9E, 16'hF75D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF5D, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hFEDD, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hDE19, 16'hE619, 16'hF69B, 16'hFE9C, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE9C, 16'hF65A, 16'hFE19, 16'hA38F, 16'hC516, 16'hFF1D, 16'hF6DD, 16'hF6DD, 16'hFF1D, 16'hFF1E, 16'hBC93, 16'hBC93, 16'hFF1D, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF71D, 16'hF6DC, 16'hEE9B,
        16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9C, 16'hEE5B, 16'hD557, 16'hEE5B, 16'hE65A, 16'hE65B, 16'hE65B, 16'hE65A, 16'hEE9B, 16'hB4D4, 16'h20C0, 16'hAD13, 16'hCDD7, 16'hC5D6, 16'hC5D6, 16'hC5D6, 16'hC5D6, 16'hC596, 16'hC5D6, 16'hC596, 16'hC5D7, 16'hCE58, 16'hCE18, 16'hD659, 16'hE69B, 16'hDE9A, 16'hBDD6, 16'hBE58, 16'hC698, 16'hBE98, 16'hC6D9, 16'h9512, 16'h8C50, 16'hE69B, 16'hEEDB, 16'h9C92, 16'hC618, 16'hE71C, 16'h734D, 16'hEEDC, 16'hC596, 16'h734D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h6B0C, 16'hE69A, 16'hE6DB, 16'hE69B, 16'hE69B, 16'hEEDC, 16'hBD55, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h8C51, 16'hAD14, 16'hB4D4, 16'hF6DC, 16'hE65A, 16'hE65A, 16'hE65A, 16'hD5D8, 16'hEE9B, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hE61A, 16'h9B4E, 16'h5B0B, 16'h83CE, 16'h30C1, 16'h93D0, 16'hE61A, 16'hFF5E, 16'hD5D7, 16'h8ACB, 16'hFE9B, 16'hFEDC, 16'hF69C, 16'hFEDD, 16'hE65A, 16'hCE9A, 16'hDF9E, 16'hCE9A, 16'hDDD8, 16'hFEDD, 16'hF69C, 16'hFEDD, 16'hFF1D, 16'hFEDD, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E,
        16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1D, 16'hFF1D, 16'hFEDD, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hFE9C, 16'hFE9C, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE9C, 16'hF65B, 16'hFE5B, 16'hDD16, 16'h938F, 16'hFEDD, 16'hF6DD, 16'hF6DD, 16'hFF1E, 16'hFEDC, 16'hB452, 16'hA38E, 16'hF69B, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DD, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hE61A, 16'hD597, 16'hEE9B, 16'hE65A, 16'hE65B, 16'hE65B, 16'hE65A, 16'hEE9B, 16'h8B8F, 16'h4A07, 16'hBD55, 16'hCDD7, 16'hC5D6, 16'hC5D6, 16'hC5D6, 16'hC5D6, 16'hC5D6, 16'hC5D6, 16'hC596, 16'hC5D6, 16'hCE18, 16'hCE18, 16'hD658, 16'hE69A, 16'hDE59, 16'h9D13, 16'hBE58, 16'hC698, 16'hBE98, 16'hC6D9, 16'h7C0F, 16'hB555, 16'hEEDB, 16'hE69B, 16'h738E, 16'hEF5D, 16'hC618,
        16'h9451, 16'hEF1C, 16'h734D, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h6B0D, 16'hDE59, 16'hEEDB, 16'hE69B, 16'hE69B, 16'hEEDC, 16'hC596, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9451, 16'hAD14, 16'hAC93, 16'hF69C, 16'hE65A, 16'hE65A, 16'hEE5B, 16'hD5D8, 16'hE65A, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC,
        16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9B, 16'hB452, 16'h4247, 16'h840F, 16'h840F, 16'h5ACA, 16'h4143, 16'h8B8E, 16'hDE18, 16'hAC51, 16'hA3D0, 16'hFEDC, 16'hFEDC, 16'hF6DC, 16'hFEDC, 16'hDE19, 16'hD659, 16'hCE18, 16'hF6DC, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hFEDD, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1D, 16'hFEDD, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hF69C, 16'hFE9C, 16'hF69B, 16'hF65B, 16'hFE9B, 16'hF65B, 16'hFE9B, 16'hF69B, 16'hF69B, 16'hFE5B, 16'hF61A, 16'h930D, 16'hE65A, 16'hFF1D, 16'hFF1D, 16'hFF1E,
        16'hDE19, 16'h9B4F, 16'hB3D0, 16'hDDD8, 16'hFEDD, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hF6DD, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hDDD9, 16'hD5D8, 16'hEE9B, 16'hE65A, 16'hE65B, 16'hE65A, 16'hEE9B, 16'hE61A, 16'h628A, 16'h6B4C, 16'hC5D6, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D6, 16'hC5D7, 16'hC5D6, 16'hC5D6, 16'hC596, 16'hAD13, 16'hCE18, 16'hCE58, 16'hCE58, 16'hDE99, 16'hCE58, 16'h8450, 16'hBE98, 16'hBE98, 16'hC698, 16'hC698, 16'h52CA, 16'hCDD7, 16'hEEDB, 16'hCE18, 16'h8410, 16'hFFDF, 16'h9492, 16'hCE18, 16'hBD96, 16'h8C10, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h734D, 16'hD619, 16'hEEDB, 16'hE69B, 16'hE69B, 16'hEEDB, 16'hCDD7, 16'h9C92, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9C92, 16'hAD13, 16'h9C11, 16'hEE9B, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hDDD8, 16'hDE19, 16'hF6DC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hF6DC, 16'hF69C, 16'hC4D5, 16'h4A07, 16'h740E, 16'h7C0E, 16'h844F, 16'h7C0F, 16'h41C7, 16'h1000, 16'hA38F, 16'h6145, 16'h938F, 16'hF65A, 16'hFEDC, 16'hFEDC, 16'hFE9C, 16'hF69B, 16'hFE9C, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hFEDD, 16'hFEDD, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hF69C, 16'hFE9C, 16'hFE9C, 16'hF65B, 16'hF69B, 16'hF65B, 16'hFE9B, 16'hF65B, 16'hFE9B, 16'hFE5A, 16'hA38F, 16'hC556, 16'hFF5E, 16'hFF1D, 16'hEE5A, 16'hB492, 16'h71C6, 16'hA34E, 16'hDD57, 16'hEE9B, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hF69C, 16'hDD98, 16'hDE19, 16'hEE9B, 16'hE65A, 16'hE65B, 16'hE65A, 16'hEE9B, 16'hCD97, 16'h3104, 16'h8C0F, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D6, 16'hC5D7, 16'hBD96, 16'h8C0F, 16'hC617, 16'hCE58, 16'hCE58, 16'hD699, 16'hC617,
        16'h740E, 16'hC698, 16'hBE98, 16'hC6D9, 16'hA594, 16'h6B4C, 16'hDE9A, 16'hEEDB, 16'hA4D3, 16'hBDD7, 16'hF79E, 16'h83CF, 16'hC5D7, 16'h5249, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h83CF, 16'hC5D7, 16'hEEDB, 16'hE69B, 16'hE69B, 16'hEEDB, 16'hD659, 16'h8410, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'hA4D3, 16'h8BD0, 16'hEE9B, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hE619,
        16'hDDD8, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF6DC, 16'hD597, 16'h5A08, 16'h6BCD, 16'h7C0F, 16'h740E, 16'h7C4F, 16'h840F, 16'h4103, 16'hDD56, 16'hE5D8, 16'h934E, 16'h828A, 16'hC4D4, 16'hE597, 16'hEE19, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hFEDD, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hF69C, 16'hFE9C, 16'hFE9C, 16'hF65B,
        16'hFE9B, 16'hF65B, 16'hFE9B, 16'hFE9B, 16'hFE5B, 16'hBC52, 16'hCD15, 16'hFE9C, 16'hDE19, 16'hB452, 16'h9B0C, 16'hCC93, 16'hABCF, 16'hBC11, 16'hE5D9, 16'hF6DD, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hD597, 16'hE65A, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hE65B, 16'hEE9B, 16'hB4D4, 16'h1840, 16'h9C91, 16'hCE17, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hB555, 16'h6B4C, 16'hC617, 16'hC658, 16'hC658, 16'hCE99, 16'hBE17, 16'h740E, 16'hC698, 16'hBE98, 16'hCED9, 16'h740E, 16'hA514, 16'hE6DB, 16'hE69B, 16'h738D, 16'hEF5C, 16'hC618, 16'h8410, 16'h5A8A, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'hB555, 16'hEEDC, 16'hE69B, 16'hE69B, 16'hE69B, 16'hDE9A, 16'h83CF, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h9451, 16'h6B0C, 16'hDE19, 16'hEE9B, 16'hE65A, 16'hE65B, 16'hE65A, 16'hD5D8, 16'hEE9B, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hF6DC, 16'hE619, 16'h728A, 16'h638C, 16'h7C4F, 16'h740F, 16'h744F, 16'h8450, 16'h3984, 16'hB493, 16'hFF1D, 16'hFE9C, 16'hEE1A, 16'hE5D8, 16'hDD97, 16'hEE19, 16'hFE9B, 16'hFE9B, 16'hFE9C, 16'hF69B, 16'hFEDC, 16'hFE9C, 16'hFEDD, 16'hF6DC, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF5E,
        16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1D, 16'hFEDD, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hFE9C, 16'hFE9C, 16'hFE9C, 16'hF69B, 16'hFE9C, 16'hFE9C, 16'hFE9B, 16'hDD97, 16'h9B4E, 16'hABD0, 16'hC493, 16'hAB8F, 16'hAB8F, 16'hCC93, 16'hED97, 16'hF5D8, 16'h9B0C, 16'hCCD4, 16'hEE5B, 16'hF6DD, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE5B, 16'hD597, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE5A, 16'h940F, 16'h4A07, 16'hA4D3, 16'hCE17, 16'hC5D7, 16'hC617,
        16'hC5D7, 16'hC5D7, 16'hC5D7, 16'hC5D6, 16'hCE17, 16'hA513, 16'h630C, 16'hC658, 16'hC658, 16'hC658, 16'hCE99, 16'hAD95, 16'h740F, 16'hC6D9, 16'hC698, 16'hBE58, 16'h52CA, 16'hCE18, 16'hE6DB, 16'hBD96, 16'h840F, 16'hF79E, 16'h7BCF, 16'h5ACB, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h9451, 16'hEEDC, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE6DB,
        16'h83CF, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8C0F, 16'h62CB, 16'hC596, 16'hEE9B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hD597, 16'hE65A, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hEEDC, 16'hEE9C, 16'hEEDC, 16'hEE9C, 16'hEEDC, 16'hF69B, 16'h938F, 16'h52CA, 16'h7C4F, 16'h744F, 16'h7C4F, 16'h8490, 16'h62CA, 16'h934E, 16'hFE9C, 16'hF65B, 16'hFE9C, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hFE9B, 16'hF65B, 16'hFE9C, 16'hF69B, 16'hFEDC, 16'hF69C, 16'hFEDD, 16'hFEDC, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hFE9C, 16'hFE9C, 16'hF65B, 16'hF65A, 16'hDD57, 16'hBC52, 16'hA34E, 16'hBC11, 16'hD4D4, 16'hD4D4, 16'hE516, 16'hED97, 16'hED97, 16'hED97, 16'hD515, 16'h8A8B, 16'hDD57, 16'hF69C, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hE619, 16'hDDD8, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hD5D8, 16'h6ACB, 16'h630B, 16'hB555, 16'hC617, 16'hC617, 16'hC617, 16'hC617, 16'hC617, 16'hC5D7, 16'hC5D6, 16'hCE18, 16'h9491, 16'h6B4D, 16'hCE98, 16'hC658, 16'hC658, 16'hCE99, 16'h9D13, 16'h8491, 16'hC6D9, 16'hC6D9, 16'h8CD2, 16'h840F, 16'hDEDB, 16'hE6DB, 16'h738D, 16'hD69A, 16'hBDD6, 16'h000, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h734D, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69A, 16'hEEDC, 16'h9C51, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h7B8E, 16'h6B0C, 16'hA493, 16'hEEDB, 16'hE65A, 16'hE65A, 16'hE65A, 16'hD5D8, 16'hDE19, 16'hEEDC, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9C, 16'hF6DC, 16'hB493, 16'h3A47, 16'h7C50, 16'h744F, 16'h7C4F, 16'h8490, 16'h738D, 16'h6A49, 16'hF65B, 16'hFE9B, 16'hF65B, 16'hF65B, 16'hF65B, 16'hF69B, 16'hFE9B,
        16'hF65B, 16'hFE9C, 16'hF69B, 16'hFEDC, 16'hFE9C, 16'hFEDD, 16'hFEDD, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFEDD, 16'hFEDD, 16'hFEDD, 16'hF69C, 16'hF69B, 16'hEE19, 16'hEE5A, 16'hFE9B, 16'hF65B, 16'hF65A, 16'hF65B, 16'hF65A, 16'hF65B, 16'hF69B, 16'hFEDD, 16'hD556, 16'h92CC, 16'hE619, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hDDD8, 16'hE619,
        16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hEE9B, 16'hA493, 16'h83CE, 16'h734D, 16'hC5D7, 16'hC617, 16'hC617, 16'hC617, 16'hC617, 16'hC617, 16'hC617, 16'hC5D7, 16'hCE18, 16'h738D, 16'h52CA, 16'hC658, 16'hC658, 16'hC658, 16'hCED9, 16'h844F, 16'h9513, 16'hCF1A, 16'hBE98, 16'h4A89, 16'hC617, 16'hE71B, 16'hBD96, 16'h8C91, 16'hD69A, 16'h000, 16'hB595, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h7BCE, 16'hCE18, 16'hEE9B, 16'hE69B, 16'hE69A, 16'hEEDB, 16'hB514, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h6B0C, 16'h734D, 16'h9C51, 16'hDE5A, 16'hE69B, 16'hE65A, 16'hE65B, 16'hDE19, 16'hD5D8, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hD597, 16'h4207, 16'h7C4F, 16'h7C50, 16'h7C90, 16'h8490, 16'h7C0F, 16'h5987, 16'hEE19, 16'hFE9B, 16'hF65A, 16'hF65B, 16'hF69B, 16'hF69B, 16'hFE9C, 16'hF69B, 16'hFEDC, 16'hF69B, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hBCD4, 16'hB410, 16'hF69B, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hDDD8, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'h7B4D, 16'h9C92, 16'h83CE, 16'hCE58, 16'hC617, 16'hC617, 16'hC617, 16'hC617, 16'hC617, 16'hC617, 16'hC617, 16'hC5D7, 16'h4A08, 16'h52CA, 16'hC658, 16'hC658, 16'hC658, 16'hC698, 16'h6BCD, 16'hAE16, 16'hCF1A, 16'h8491, 16'h8C51, 16'hDEDA, 16'hDEDA, 16'h7BCE, 16'h9D13, 16'h31C6, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'hA493, 16'hEEDC, 16'hE69A, 16'hE69B, 16'hE6DB, 16'hCE18, 16'h8C51, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9492, 16'h6ACB, 16'h9C92, 16'hBD56, 16'hEE9B, 16'hE65A, 16'hE65B, 16'hE65A, 16'hCD97, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF69C, 16'hEE5A, 16'h628A, 16'h740E,
        16'h8490, 16'h7C90, 16'h8490, 16'h8490, 16'h49C6, 16'hE619, 16'hFE9C, 16'hF65A, 16'hFE9B, 16'hF69B, 16'hF69B, 16'hFE9C, 16'hF69B, 16'hFEDC, 16'hFEDC, 16'hFEDC, 16'hFEDD, 16'hFEDD, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF1E, 16'hFF5E, 16'hFF1D, 16'h8B4D, 16'hCD56, 16'hF6DC, 16'hF6DC, 16'hF6DC, 16'hEEDC, 16'hEE9B, 16'hEE9B, 16'hEE9B,
        16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5A, 16'hDE19, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hEE9B, 16'hB4D4, 16'h8C10, 16'h9C92, 16'h9491, 16'hCE58, 16'hC617, 16'hC617, 16'hC617, 16'hC617, 16'hC617, 16'hC617, 16'hC617, 16'hB595, 16'h3186, 16'h634C, 16'hC658, 16'hC698, 16'hC698, 16'hB616, 16'h530A, 16'hC6D9, 16'hADD6, 16'h4A89, 16'hCE59, 16'hE71C, 16'h9CD3, 16'h080, 16'h6B4C, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h6B0C, 16'hE69B, 16'hE69A, 16'hE69B, 16'hE69A, 16'hE69A, 16'h83CF, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h41C7, 16'hBD95, 16'h8BD0, 16'hEE9B, 16'hE65A, 16'hE65A, 16'hE65A, 16'hD597, 16'hDE19, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF69C, 16'h8BCF, 16'h5B4C, 16'h84D1, 16'h7C90, 16'h8490, 16'h8CD1, 16'h4206, 16'hCD57, 16'hFEDD, 16'hF65A, 16'hFE9C, 16'hF69B, 16'hF69B, 16'hFE9C, 16'hFEDC, 16'hFEDC, 16'hFEDD, 16'hFEDD, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E,
        16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hD5D7, 16'h6986, 16'hE619, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hE65A, 16'hEE9B, 16'h730C, 16'hBD55, 16'h8C10, 16'hAD54, 16'hCE58, 16'hC617, 16'hC617, 16'hC617, 16'hC617, 16'hC617, 16'hC617, 16'hCE58, 16'h9CD2, 16'h7C0F, 16'h7BCF, 16'hBE58, 16'hC698, 16'hCED9, 16'h9D54, 16'h7C0F, 16'hCED9, 16'h4248, 16'hAD55, 16'hE71C, 16'h9D13, 16'h31C6, 16'hC617, 16'hF79E,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h8410, 16'hBD96, 16'hEEDB, 16'hE69A, 16'hE69A, 16'hEEDB, 16'h9451, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h000, 16'hCE18, 16'h7B8E, 16'hDE19, 16'hEE9B, 16'hE65A, 16'hEE9B, 16'hDDD8, 16'hD5D7, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B,
        16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF6DC, 16'hBD14, 16'h3A88, 16'h84D1, 16'h8491, 16'h8491, 16'h8CD2, 16'h4A88, 16'hC515, 16'hFF1D, 16'hF69B, 16'hFEDC, 16'hF6DC, 16'hFEDC, 16'hFEDC, 16'hFEDD, 16'hFEDD, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E,
        16'hFF5E, 16'hFF1D, 16'h7289, 16'h9B8E, 16'hF69B, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hE65A, 16'hE65B, 16'hE65B, 16'hE65A, 16'hEE9B, 16'hBD55, 16'h7B4E, 16'hCDD7, 16'h630B, 16'hC617, 16'hC657, 16'hC657, 16'hC617, 16'hC617, 16'hC617, 16'hC617, 16'hC617, 16'hCE58, 16'h738D, 16'hBE17, 16'h8C50, 16'hBE57, 16'hCE99, 16'hCED9, 16'h73CE, 16'h9D13, 16'h8450, 16'h9CD2, 16'hD6DA, 16'h738D, 16'h5289, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h62CB, 16'hE69B, 16'hE69A, 16'hE69A, 16'hEEDB, 16'hBD96, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h5ACB, 16'hBDD6, 16'h840F, 16'hACD3, 16'hEE9C, 16'hE65A, 16'hEE5B, 16'hE619, 16'hCD96, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hF6DC, 16'hDE19, 16'h4247, 16'h84D1, 16'h84D1, 16'h84D1, 16'h8D12, 16'h5B0B, 16'hA411, 16'hFF1D, 16'hFEDD, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E,
        16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hC515, 16'h000, 16'hCD15, 16'hF6DC, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hE65A, 16'hE65A, 16'hE65B, 16'hE65B, 16'hE65A, 16'hEE9B, 16'h72CC, 16'hC556, 16'hBD55, 16'h7BCF, 16'hCE58, 16'hC617, 16'hC657, 16'hC617, 16'hC617, 16'hC617, 16'hC617, 16'hC617, 16'hC617, 16'h630C, 16'hDEDB, 16'h7BCE, 16'hBE57,
        16'hCED9, 16'hC658, 16'h52CA, 16'h5B0B, 16'h6BCD, 16'h9D13, 16'h5ACA, 16'h9D13, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9451, 16'hAD14, 16'hEEDB, 16'hDE9A, 16'hE69B, 16'hDE5A, 16'h734D, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'h9CD2, 16'hA513,
        16'hAD55, 16'h4208, 16'hE69A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hCD96, 16'hDE19, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9C, 16'hF69C, 16'hEE9B, 16'h6B0C, 16'h744F, 16'h8D12, 16'h84D1, 16'h84D2, 16'h740E, 16'h728A, 16'hF6DC, 16'hFF1E, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1D, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E,
        16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hE65A, 16'h5000, 16'h6A08, 16'hE61A, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hE65A, 16'hE65B, 16'hE65B, 16'hE65A, 16'hEE9B, 16'hB515, 16'h7B4D, 16'hE659, 16'h8C0F, 16'hAD55, 16'hC658, 16'hC617, 16'hC617, 16'hC657, 16'hC657, 16'hC617, 16'hC617, 16'hCE58, 16'hA554, 16'h8410, 16'hFFDF, 16'h73CE, 16'hBE57, 16'hD6DA, 16'hAD95, 16'h000, 16'h4A89, 16'h8C91, 16'hB596, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h4A08, 16'hD618, 16'hE6DB, 16'hDE9A, 16'hEEDB, 16'hA493, 16'hBD97, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h83CF, 16'hCE18, 16'h000, 16'hB555, 16'hEE9B, 16'hE65A, 16'hEE9B, 16'hDE18, 16'hCD96, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE9C, 16'hEE9B, 16'hF6DC, 16'hA492, 16'h538C, 16'h8D12, 16'h84D1, 16'h84D2, 16'h8CD2, 16'h4144, 16'hDE19, 16'hFF5F, 16'hFF1E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E,
        16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hF71C, 16'h7A8A, 16'h4183, 16'h9C10, 16'hF69C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hE65A, 16'hE65B, 16'hE65A, 16'hE65B, 16'hDE19, 16'h5A09, 16'hC596, 16'hD618, 16'h7B8E, 16'hC618, 16'hC658,
        16'hC658, 16'hC657, 16'hC657, 16'hC657, 16'hC657, 16'hC617, 16'hCE98, 16'h7BCE, 16'hBDD7, 16'hFFDF, 16'h7BCF, 16'hBE57, 16'hD71A, 16'h73CE, 16'hB596, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hD65A, 16'h628A, 16'hDE9A, 16'hE69B, 16'hE69B, 16'hDE5A, 16'h6B0C, 16'hEF5D, 16'hFFDF, 16'hF79E, 16'h738D, 16'hC5D7, 16'h5B4C, 16'h4ACA, 16'hD618, 16'hEE9B, 16'hE65A, 16'hE65A, 16'hC555, 16'hE65A, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hEE9C, 16'hEE9B, 16'hF6DC, 16'hCD97, 16'h4AC9, 16'h8D12, 16'h84D2, 16'h84D2, 16'h8D12, 16'h52C9, 16'hAC93, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hF71D, 16'hF71D, 16'hFF1D, 16'hF71D, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF5E, 16'h9BCF, 16'h630B, 16'h5A89, 16'hCD56, 16'hF69C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hE65A, 16'hE65A, 16'hE65B, 16'hE65A, 16'hEE9B, 16'h9C11, 16'h730C, 16'hE69A, 16'hACD3, 16'h9CD2, 16'hCE98, 16'hC657, 16'hC658, 16'hC658, 16'hC657, 16'hC657, 16'hC657, 16'hC658, 16'hBE17, 16'h634C, 16'hEF9D, 16'hFFDF, 16'h8410, 16'hC698, 16'hC698, 16'h73CE, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h734D, 16'hE6DB, 16'hE69B, 16'hEEDB, 16'hA4D3, 16'hB556, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h9450, 16'h7C50, 16'h5C4E, 16'h6B4D, 16'hE65B, 16'hEE5B, 16'hEE9B, 16'hCD97, 16'hD5D7, 16'hEE9B, 16'hE69A, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hEE9B, 16'hEE9B, 16'hEE9C, 16'hEE5B, 16'h6B0B, 16'h7C90, 16'h8D12, 16'h84D2, 16'h8D12, 16'h8491, 16'h6A48, 16'hF6DC,
        16'hFF5F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hDE19, 16'hDDD8, 16'hF6DC, 16'hFEDC, 16'hEE5A, 16'hDDD8, 16'hF71C, 16'hFF9F, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hAC52, 16'h5206, 16'h8C90, 16'h6249, 16'hEE5A, 16'hEE9C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A,
        16'hE65A, 16'hE69A, 16'hE65A, 16'hEE9B, 16'hCDD7, 16'h000, 16'hB555, 16'hDE9A, 16'h8C50, 16'hBE17, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hBE57, 16'hCE98, 16'h9491, 16'h94D2, 16'hFFDF, 16'hF79E, 16'h73CE, 16'hCE99, 16'h8C91, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h730C, 16'hD659, 16'hEEDB, 16'hE69A, 16'h6B4C, 16'hDEDB, 16'hFFDF, 16'hDEDB, 16'h5ACA, 16'h6B8D, 16'h9E15, 16'h5C4E, 16'h9C51, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hC556, 16'hE69A, 16'hE69B, 16'hE65B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hE65B, 16'hE65B, 16'hEE9B, 16'hEE9B, 16'hF6DC, 16'hA492, 16'h5B8C, 16'h8D13, 16'h84D2, 16'h8512, 16'h9553, 16'h5ACA, 16'hB4D4, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hF71D, 16'hD618, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF71D, 16'hDE19, 16'hFF5E, 16'hFF9F,
        16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF9F, 16'hB493, 16'h3800, 16'h9D53, 16'h6B8D, 16'h9B8F, 16'hF69C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hE65A, 16'hE61A, 16'hE65A, 16'hE65A, 16'hE69B, 16'hE65A, 16'h628B, 16'h3185, 16'hDE59, 16'hC5D6, 16'hA554, 16'hCE99, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hBE58, 16'hC658, 16'h52CA, 16'hDEDA, 16'hFFDF, 16'hE71C, 16'h634C, 16'hB5D6, 16'h6B8E, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE18, 16'h630C, 16'hBD95, 16'hEF1C, 16'hCDD7, 16'h62CB, 16'hF75E, 16'hFFDF, 16'h8410, 16'h000, 16'h9E15, 16'hB6D8, 16'h2A06, 16'hC556, 16'hEE9B, 16'hEE9B, 16'hCD96, 16'hD5D8, 16'hEE9B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE65B, 16'hE65B,
        16'hE65B, 16'hE65B, 16'hEE9B, 16'hF69C, 16'hCDD8, 16'h4AC9, 16'h8D12, 16'h8D12, 16'h8D12, 16'h8D12, 16'h8D12, 16'h5A46, 16'hE659, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF9E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF5E, 16'hAC52, 16'h4100, 16'h9D53, 16'hA594, 16'h5A48, 16'hCD56, 16'hF69C, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B,
        16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hD5D8, 16'hDE1A, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hACD3, 16'h000, 16'h9451, 16'hDE9A, 16'hAD54, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hBE57, 16'hC699, 16'h94D2, 16'h73CE, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h6B8D, 16'h638D, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h9451, 16'h9C92, 16'hC5D7, 16'hAD14, 16'h8C10, 16'hFFDF, 16'hDF1B, 16'h000, 16'h7490, 16'hBF1A, 16'h6C4F, 16'h6A4A, 16'hEE5A, 16'hEE9B, 16'hE659, 16'hC556, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69B, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'h738D, 16'h7490, 16'h8D53, 16'h8D12, 16'h8D12, 16'h8D53, 16'h8491, 16'h6208, 16'hEEDB, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hF71C, 16'h934E, 16'h6287, 16'hADD5, 16'hAE16, 16'h8CD1, 16'h728A, 16'hEE5A, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hDE19, 16'hCD96, 16'hEE9B, 16'hE65A, 16'hEE9B, 16'hD5D8, 16'h41C7, 16'h31C6, 16'hBDD6, 16'hD659, 16'hBE17, 16'hC698, 16'hBE57, 16'hC658, 16'hC658, 16'hC658, 16'hC658, 16'hBE57, 16'hC658, 16'hB5D7, 16'h000, 16'hD699, 16'hFFDF, 16'hFFDF, 16'h8C91, 16'h000, 16'h9D13, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hE71C, 16'hD69A, 16'hCE59, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h9CD2, 16'h9CD2, 16'h6B4C, 16'h7B8E, 16'hE71C, 16'h9492, 16'h182, 16'hAE98, 16'h9E15, 16'h000, 16'h9C92, 16'hEEDB,
        16'hEE9B, 16'hCD96, 16'hD5D7, 16'hE69B, 16'hE69A, 16'hE69A, 16'hE69B, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hF69C, 16'hB514, 16'h4B4B, 16'h9553, 16'h8D13, 16'h8D53, 16'h8D12, 16'h9594, 16'h8490, 16'h6A08, 16'hE69A, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hDE19, 16'h6A08, 16'h7C0E,
        16'hB616, 16'hAE56, 16'hA5D5, 16'h6B8C, 16'hB492, 16'hF69B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65B, 16'hEE9B, 16'hB4D4, 16'hDDD8, 16'hEE9B, 16'hE65A, 16'hEE9B, 16'h9410, 16'h4A89, 16'h738D, 16'hD699, 16'hCE99, 16'hCED9, 16'hB616, 16'hADD5, 16'hC698, 16'hC658, 16'hC658, 16'hBE57, 16'hC698, 16'hB616, 16'h4248, 16'h6B8D, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h000, 16'h8450, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hEF5D, 16'hD6DB, 16'hC618, 16'hB596, 16'hA514, 16'h9492, 16'h8C51, 16'h8C51, 16'h8410, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hD69A, 16'hBDD7, 16'hBDD7, 16'hD69A, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hC618, 16'h8C50, 16'h3185, 16'h73CE, 16'h000, 16'h7CD0, 16'hBF19, 16'h6C0E, 16'h3A48, 16'hBD15, 16'hF6DC, 16'hDE59, 16'hBD14, 16'hE65A, 16'hE69B, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hDE59, 16'h4A89, 16'h8512, 16'h8D53, 16'h8D53, 16'h8D53, 16'h8D53, 16'h9DD5, 16'h8491, 16'h4901, 16'hD5D7, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E,
        16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hF6DC, 16'hAC11, 16'h6186, 16'hA553, 16'hB697, 16'hAE56, 16'hAE16, 16'h9D93, 16'h6289, 16'hDDD8, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'hCD97, 16'hA452, 16'hEE9B, 16'hE65A, 16'hEE9B, 16'hCD97, 16'h5B0B, 16'h840F, 16'hA513, 16'hDEDA, 16'hCEDA, 16'hC699, 16'h840F, 16'hB616, 16'hC698, 16'hC658, 16'hBE58, 16'hCE99, 16'hADD5, 16'h7C0F, 16'h5B0B, 16'hCE59, 16'hFFDF, 16'hEF9D,
        16'h8C1, 16'h8C50, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hAD55, 16'h9CD3, 16'h8C51, 16'h8410, 16'h8410, 16'h8C51, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'h8410, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h9492, 16'h8410, 16'h8C51, 16'h8C51, 16'h8410, 16'h9CD3, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hC618, 16'h8C51, 16'h000, 16'h9D94, 16'h8D12, 16'h94D2, 16'h6B8D, 16'hD5D8, 16'hEEDB, 16'hD5D7, 16'hCD97, 16'hE69B, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hEE9B, 16'h9411, 16'h538C, 16'h9594, 16'h8D53, 16'h8D53, 16'h8D53, 16'h9594, 16'h9DD5, 16'h8D12, 16'h2901, 16'hA451, 16'hF71D, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hCD56, 16'h7A49, 16'h840E, 16'hB656, 16'hB697, 16'hAE56, 16'hAE56, 16'hAE56, 16'h740E, 16'hA451, 16'hEE9B, 16'hE65B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hEE9B, 16'h93CF, 16'hD5D8, 16'hEE9B, 16'hE65A, 16'hEE9B, 16'h7B8E, 16'hB595, 16'h6B8D, 16'hCE58, 16'hE71B, 16'hCE99, 16'h7C0F, 16'h7C0F, 16'hCE98, 16'hC658, 16'hC698, 16'hCED9, 16'hA554, 16'h6B8D, 16'hA514, 16'h8410, 16'hFFDF, 16'hF79E, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h8410, 16'h9492, 16'h9492, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h9CD3,
        16'hAD55, 16'hC618, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'hCE59, 16'hCE59, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h8C51, 16'h9492, 16'h8C51, 16'h8C51, 16'h9492, 16'h8C51, 16'h9CD3, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF7DE, 16'h634C, 16'h52CA, 16'h4AC9, 16'h73CE, 16'h8C91, 16'h6ACB, 16'hCD97, 16'hD618, 16'hCDD7, 16'hDE59, 16'hE69A, 16'hE69A, 16'hE69A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hCDD8, 16'h19C3, 16'h8512, 16'h9594, 16'h8D93, 16'h9593, 16'h9594, 16'h95D4, 16'hA5D5, 16'h9D94, 16'h5B4B, 16'h6A49, 16'hC596, 16'hFF5E,
        16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hD5D7, 16'h8B0C, 16'h7B4B, 16'hAE15, 16'hBED8, 16'hB697, 16'hAE56, 16'hAE56, 16'hAE56, 16'h9DD4, 16'h730B, 16'hE619, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5A, 16'hF69B, 16'hB4D4, 16'h8BCF, 16'hEE9B, 16'hE65A, 16'hEEDB, 16'hACD3, 16'h9CD3, 16'hCE58, 16'h94D2, 16'hDF1B, 16'hA554, 16'h7BCE, 16'h4A88,
        16'hAD95, 16'hCE99, 16'hCE99, 16'hC698, 16'h7C4F, 16'h73CE, 16'hDF1B, 16'h6B4D, 16'hD69A, 16'hFFDF, 16'hE71C, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8C51, 16'h8C51, 16'h9492, 16'hA514, 16'h9CD3, 16'h9492, 16'h8C51, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h9CD3, 16'h8410, 16'h8C51, 16'h8410, 16'h8410, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8C51, 16'h9492, 16'h8C51, 16'hC618, 16'hC618, 16'h8C51, 16'h9492, 16'h8410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h7C50, 16'hB596, 16'h2A06, 16'hBDD7, 16'h7BCF, 16'hB514, 16'hDE18, 16'hDE19, 16'hDE59, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hEE9B, 16'h7B8E, 16'h430A, 16'h9594, 16'h9594, 16'h9594, 16'h9594, 16'h9DD4, 16'h9DD4, 16'h9DD5, 16'hA615, 16'h8D13, 16'h5289, 16'h7B0C, 16'hD5D8, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hD5D8, 16'h934D, 16'h72CA, 16'hA593, 16'hC6D8, 16'hBED8, 16'hB697, 16'hB697, 16'hB697, 16'hAE56, 16'hB696, 16'h7C4E, 16'hBCD4, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hE65A, 16'hEE9B, 16'hDDD8, 16'h3083, 16'hCD97, 16'hE69A, 16'hE69A, 16'hDE59, 16'h5A89, 16'hE75C, 16'h8410, 16'h8C51, 16'h7BCF, 16'h9491, 16'h7BCE, 16'h8C91, 16'hD6DA, 16'hC658, 16'h9D12, 16'h5B0B, 16'hAD95, 16'hF79E, 16'h8410, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hEF5D, 16'hF79E, 16'hFFDF, 16'hBDD7, 16'h8C51, 16'h8C51, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h8C51, 16'h9492, 16'h8C51, 16'h8C51, 16'h9492, 16'h8410, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h8C51, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8C51, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h7C0F, 16'hBE18, 16'h9D13, 16'hC618, 16'hEF5D, 16'h838E, 16'hE659, 16'hDE59, 16'hB514, 16'hE65A, 16'hE69A, 16'hE65A, 16'hE65A, 16'hE69A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hBD96,
        16'h0C0, 16'h7CD0, 16'h9DD4, 16'h9593, 16'h9594, 16'h9DD5, 16'h9DD5, 16'h9DD5, 16'h9DD5, 16'hA615, 16'hA615, 16'h84D1, 16'h52C9, 16'h8B4D, 16'hD5D8, 16'hF75D, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hD597, 16'h8ACC, 16'h7B0B, 16'hA593, 16'hC6D8, 16'hC718, 16'hBED7, 16'hB696, 16'hB697, 16'hB697, 16'hAE56, 16'hB697, 16'h9DD3, 16'hA410, 16'hE619, 16'hE65A, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hEE5B, 16'hE65A, 16'hEE9B, 16'hE659, 16'h5A09, 16'h7B4D,
        16'hDE5A, 16'hE65A, 16'hEEDB, 16'h7B8E, 16'hC618, 16'hE71C, 16'h630B, 16'hAD95, 16'hD699, 16'hAD95, 16'h738D, 16'hB595, 16'h8C50, 16'h634C, 16'hA514, 16'hEF5D, 16'hFFDF, 16'h7BCF, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h8C51, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h8C51, 16'h9492, 16'h8C51, 16'hBDD7, 16'hAD55, 16'h8C51, 16'h9492, 16'h8410, 16'hE71C, 16'hFFDF, 16'hCE59, 16'h8C51, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h5B4B, 16'hC658, 16'h52CA, 16'hF79E, 16'hD69A, 16'h8BD0, 16'hE69B, 16'h9C92, 16'h9C92, 16'hE6DB, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'h6B4C, 16'h2A06, 16'h8512, 16'h9DD4, 16'h9594, 16'h9DD5, 16'h9DD5, 16'h9DD5, 16'h9DD5, 16'h9DD5, 16'hA615, 16'hAE56, 16'hAE56, 16'h8D12, 16'h5288, 16'h7A89, 16'hC556, 16'hEEDC, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hD597, 16'h8B0C, 16'h7ACA, 16'hAD93, 16'hC6D8, 16'hC718, 16'hBED8, 16'hBED7, 16'hBED7, 16'hA614, 16'hB697, 16'hB697, 16'hB697, 16'hAE56, 16'h9450, 16'hDD98, 16'hD597, 16'hEE5A, 16'hEE5B, 16'hEE9B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hE65B, 16'hEE5B, 16'hEE9B, 16'hEE9B, 16'hEE9B, 16'hE65A, 16'hEE9B, 16'hDE19, 16'h72CC, 16'h1000, 16'hCDD7, 16'hE69A, 16'hEEDC, 16'hB555, 16'h840F, 16'hFFDF, 16'hAD55, 16'hE71C, 16'hFFDF, 16'hC617, 16'h4A49, 16'h9CD2, 16'h9CD2, 16'hBDD7, 16'hF79E, 16'hFFDF, 16'hDEDB, 16'h7BCF, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h8C51, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8C51, 16'h8C51, 16'hC618, 16'hFFDF, 16'hBDD7, 16'h8C51, 16'h8410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h7C0F, 16'h9D13, 16'hAD55, 16'hFFDF, 16'hAD14, 16'hA493, 16'hD618, 16'h1900, 16'h9C92, 16'hE69A,
        16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hB514, 16'h638C, 16'h5B8C, 16'h8552, 16'h9E15, 16'h9DD4, 16'h9E15, 16'h9E15, 16'h9E15, 16'h9DD5, 16'h9594, 16'hA616, 16'hA656, 16'hAE97, 16'hB657, 16'h9D53, 16'h3080, 16'h6A07, 16'h9C10, 16'hDE59, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hF71D, 16'hC596, 16'h72CB, 16'h734B, 16'hADD4, 16'hC6D8, 16'hC6D8, 16'hBED8, 16'hBED8, 16'hBED8, 16'hBED8, 16'hB696, 16'h9DD3, 16'hBED7, 16'hB697, 16'hB697, 16'h9490, 16'hD597, 16'hCD15, 16'hDDD8, 16'hEE9B, 16'hE65A, 16'hEE9B, 16'hEE5B, 16'hEE5B,
        16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE9B, 16'hE65A, 16'hEE5B, 16'hF69C, 16'hCD97, 16'h730C, 16'h4186, 16'h838E, 16'hE659, 16'hEEDB, 16'hD619, 16'h4A08, 16'hEF5D, 16'hF79E, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hEF9D, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hCE59, 16'hC618, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF9E, 16'h9492, 16'h9492, 16'h9492, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8C51, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8C51, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hBDD7, 16'h8C51, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h9CD3, 16'hF7DF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h73CE, 16'h7C0F, 16'h8CD1, 16'hEF5D, 16'hFFDF, 16'h6B0C, 16'hC596, 16'hA492, 16'h5AC9, 16'h8C10, 16'hE65A, 16'hE69A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hD619, 16'h73CE, 16'hB617, 16'h4B0A, 16'h8D93, 16'hA615, 16'h9E15, 16'h9E15, 16'hA656, 16'h9593, 16'h7CD1, 16'hAE57, 16'hA656, 16'hAE56, 16'hB697, 16'hAE56, 16'h8450, 16'hA513, 16'h5B0A, 16'h6A89, 16'h82CB, 16'hBD15, 16'hEEDC, 16'hFF5E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hE69B, 16'hACD3, 16'h49C7, 16'h000, 16'h000, 16'hA5D4, 16'hCF59, 16'hC718, 16'hA593, 16'hB656, 16'hBED8, 16'hBED7, 16'hC6D8, 16'h9D92, 16'hB656, 16'hBED8, 16'hB697, 16'h9CD1, 16'hBC93, 16'hBC93, 16'hB493, 16'hEE5B, 16'hEE5A, 16'hEE5A, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hEE5B, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hEE9B, 16'hA452, 16'h6B0C, 16'hBD56, 16'h49C7, 16'hCD96, 16'hEEDB, 16'hE6DB, 16'h5A49, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h9492, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8C51, 16'h8C51, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h8C51, 16'hA514, 16'hFFDF, 16'hC618, 16'h8C51, 16'h8C51, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8C51, 16'h8C51, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hF79E, 16'h8450, 16'h11C2, 16'hB5D6, 16'hFFDF, 16'hD6DA, 16'h6B0C, 16'hC5D6, 16'hAD14, 16'hB596, 16'h738D, 16'hDE5A, 16'hE65A, 16'hDE5A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hA4D3, 16'hA554, 16'hDEDB, 16'h1204, 16'h9593, 16'hA656, 16'h9E15, 16'hAE57, 16'h9553, 16'h4309, 16'hAE56, 16'hAE56, 16'hAE56, 16'hAE97, 16'hB697, 16'h7C50, 16'hCE99, 16'h7C90, 16'hBE98, 16'hA594, 16'h7BCE, 16'h6A88, 16'h938D, 16'hBD14, 16'hE69A, 16'hFF5E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFFDF, 16'hFF5E, 16'hD619, 16'h8C10, 16'h000, 16'h000, 16'h000, 16'h2104, 16'h000, 16'hADD5, 16'hC718, 16'hC718, 16'h94D0, 16'hADD5, 16'hCF19, 16'hA5D4, 16'h94D1, 16'hA512, 16'hBE16,
        16'hADD5, 16'h9C90, 16'hAC10, 16'h934E, 16'h724A, 16'hE65A, 16'hEE9B, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5B, 16'hE65A, 16'hE65B, 16'hEE9B, 16'hEE9B, 16'hCD96, 16'h72CC, 16'hA493, 16'hEF1C, 16'h734D, 16'h9410, 16'hEEDB, 16'hE69B, 16'h7B4D, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8C51, 16'h8410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8C51, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hDEDB, 16'h8C51, 16'h8C51, 16'hA514, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h8C51, 16'hD69A, 16'hF79E, 16'hCE59, 16'h8C51, 16'h9492, 16'h8410, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD95, 16'h1983, 16'hD69A, 16'hFFDF, 16'hBDD7, 16'h7BCF, 16'h8C91, 16'hDEDB, 16'hCE59, 16'h5A89, 16'hD618, 16'hE69A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE69A, 16'h634B, 16'hD6DB, 16'hDF1B, 16'h203, 16'h9DD5, 16'hAE97, 16'hAE57, 16'h9D94, 16'h63CD, 16'h84D1, 16'hB697, 16'hAE57, 16'hB697, 16'hBED8, 16'h6C0E, 16'hE71C, 16'hA554, 16'h9593,
        16'hCF5A, 16'hC719, 16'hBE98, 16'hA594, 16'h738C, 16'h6AC9, 16'h8B4C, 16'hAC92, 16'hD618, 16'hF71C, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hE6DB, 16'hB555, 16'h62CB, 16'h000, 16'h000, 16'h041, 16'h20C4, 16'h1082, 16'h000, 16'h20C3, 16'hB657, 16'hC718, 16'hC718, 16'h840E, 16'h9491, 16'hBED7, 16'hCF18, 16'h840E, 16'h6ACA, 16'h6247, 16'h3800, 16'h834D, 16'hCDD7, 16'h624A, 16'hC556, 16'hEE9B, 16'hE65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hE65A, 16'hE65A, 16'hEE9B, 16'hEE5A, 16'hCD97, 16'h8B8F, 16'h3985, 16'hDE99, 16'hFF9E, 16'h7BCF, 16'h6B0C, 16'hEF1B, 16'hDE9A, 16'h6ACB, 16'hAD54, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8C51, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8C51, 16'h8C51, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8C51, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h8C51, 16'h9492, 16'h8C51, 16'h9492, 16'h8C51, 16'h9492, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDF1B, 16'h8450, 16'hC658, 16'hFFDF, 16'hB595, 16'h5B0A, 16'h738E, 16'hFFDF, 16'hCE59, 16'h5248, 16'hC5D7, 16'hDE59, 16'hE69A, 16'hE65A, 16'hDE59, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE65A, 16'hE659, 16'hE69A, 16'hCDD8, 16'h530A, 16'hFFDF, 16'hD69A, 16'h2246, 16'hAE16, 16'hBED9, 16'h8512, 16'hC659, 16'h9D54, 16'h8D52, 16'hBED8, 16'hAE57, 16'hC6D9, 16'h748F, 16'hCE59, 16'hF7DF, 16'h5B8C, 16'hBE98, 16'hC719, 16'hC719, 16'hC71A, 16'hCF19, 16'hC6D9, 16'hB616, 16'h94D1, 16'h3983, 16'h6ACA, 16'h9C50, 16'hBD14, 16'hDE19, 16'hFF5D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF71D, 16'hCDD8, 16'h83CF, 16'h000, 16'h000, 16'h000, 16'h18C3, 16'h18C3, 16'h800, 16'h000, 16'h000,
        16'h000, 16'h1040, 16'hBE16, 16'hCF1A, 16'hCF5A, 16'h9CD1, 16'h8C50, 16'h9D53, 16'h8CD0, 16'h948F, 16'h9490, 16'hAD14, 16'hD699, 16'hF75D, 16'h9451, 16'hAC93, 16'hF69B, 16'hE65A, 16'hEE5A, 16'hEE5A, 16'hEE5A, 16'hEE5B, 16'hF69B, 16'hEE9B, 16'hC555, 16'hA451, 16'h838D, 16'h83CF, 16'hFF9E, 16'hF75D, 16'h5ACA, 16'h8C10, 16'hEEDB, 16'hBD96, 16'h62CA, 16'hC5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hD69A, 16'h8410, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8410, 16'h9492, 16'h9492, 16'hE71C, 16'hFFDF, 16'hCE59, 16'h8C51, 16'h9492, 16'h8410, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h9492, 16'h8410, 16'h9492, 16'h9492, 16'h9492, 16'h8410, 16'h9CD3, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'hE71B, 16'hFFDF, 16'hC617, 16'h2942, 16'h9491, 16'hFFDF, 16'hD699, 16'h630A, 16'h9C91, 16'hB514, 16'hDE19, 16'hE69A, 16'hE65A, 16'hE659, 16'hE659, 16'hE659, 16'hE659, 16'hDE59, 16'hE69B, 16'hAD14, 16'h8C90, 16'hFFDF, 16'hCE99, 16'h3A88,
        16'hBE98, 16'h9DD4, 16'hBE18, 16'hFFDF, 16'h7C0F, 16'h9593, 16'hBED8, 16'hC719, 16'h9593, 16'h9D14, 16'hFFDF, 16'hC658, 16'h5BCC, 16'hC719, 16'hC6D9, 16'hBED8, 16'hBED9, 16'hC719, 16'hCF5A, 16'hD79B, 16'hBE57, 16'h73CE, 16'h8C50, 16'h6B0A, 16'h83CE, 16'h6A49, 16'h938F, 16'hBD55, 16'hEEDC, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF5E, 16'hDE5A, 16'hA4D3, 16'h41C7, 16'h000, 16'h000, 16'h000, 16'h2104, 16'h1082, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h041, 16'h000, 16'h6B4C, 16'hB5D5, 16'hBE57, 16'h9C91, 16'h840F, 16'hF79D, 16'hBD55, 16'hBD95, 16'hD658, 16'hEF1C, 16'hCE59, 16'h7B8E, 16'hAC93, 16'hEE5B, 16'hE65A, 16'hEE5A, 16'hEE9B, 16'hF69B, 16'hF69B, 16'hE619, 16'hC514, 16'h8B8E, 16'hAD14, 16'hDE9A, 16'h9C92, 16'hEF1C, 16'hD659, 16'h4A08, 16'h9C91, 16'hBD55, 16'h8C10, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h9CD3, 16'hF79E, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h9CD3, 16'h8C51, 16'h9492, 16'h8410, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hB596, 16'h9492, 16'h8C51, 16'h9492, 16'hBDD7, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h4A49, 16'h9491, 16'hFFDF, 16'hDEDB, 16'h738D, 16'h8410, 16'h8C10, 16'hA493, 16'hD618, 16'hE69A, 16'hE69A, 16'hE659, 16'hDE59, 16'hDE19, 16'hDE19, 16'hE69A, 16'hAD13, 16'h9D13, 16'hFFDF, 16'hD6DA, 16'h740E, 16'h84D1, 16'hA554, 16'hFFDF, 16'hF79E, 16'h8450, 16'h84D1, 16'hBED8, 16'hC6D9, 16'h7C50, 16'hF79E, 16'hFFDF, 16'hAD96, 16'h5BCC, 16'hC6D9, 16'hC71A, 16'hC719, 16'hC719, 16'hCF1A, 16'hCF1A, 16'hDF9C, 16'hCED9, 16'h94D1, 16'h8C90, 16'hE71B, 16'hDEDB, 16'hAD95, 16'h5ACA, 16'h800, 16'h5A08, 16'h9410, 16'hC556, 16'hEE9B, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hE69A, 16'hB555, 16'h6B0C, 16'h000,
        16'h000, 16'h000, 16'h18C3, 16'h18C3, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h5A89, 16'h734C, 16'h4A07, 16'h62CA, 16'h6B0B, 16'h6B0B, 16'hB554, 16'hACD3, 16'h834D, 16'h59C7, 16'h834D, 16'hD5D8, 16'hFEDC, 16'hF69B, 16'hF6DC, 16'hEE5A, 16'hDDD8, 16'hC515, 16'hAC51, 16'h8B8E, 16'hAD14, 16'hEF5C, 16'hEF5C, 16'h7B8D, 16'h6B0B, 16'hAD14, 16'hAD14, 16'hCE18, 16'hBD96, 16'hA4D3, 16'hDEDA, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h8410, 16'h9CD3, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hEF5D, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9CD2, 16'hA514, 16'hFFDF, 16'hEF5D, 16'h9CD3, 16'h840F, 16'h7BCE,
        16'h630B, 16'h9410, 16'hC596, 16'hDE59, 16'hE69A, 16'hE69A, 16'hE65A, 16'hDE59, 16'hE6DA, 16'hAD54, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hA555, 16'h8C91, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD96, 16'h63CD, 16'h8D12, 16'h4B0A, 16'hB5D7, 16'hFFDF, 16'hFFDF, 16'hAD95, 16'h534A, 16'hAE16, 16'hCF1A, 16'hCF1A, 16'hCF1A, 16'hC6D9, 16'hBE57, 16'hADD5, 16'hAD94, 16'h5A48, 16'h800, 16'h840F, 16'h8C50, 16'h7B8D, 16'h62CA, 16'h83CE, 16'h840F, 16'h6B0A, 16'h5904, 16'h8B0D, 16'hC555, 16'hE659, 16'hE65A, 16'hD618, 16'hB515, 16'h7B8E, 16'h000, 16'h000, 16'h000, 16'h18C3, 16'h20C3, 16'h841, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h841, 16'h000, 16'h2144, 16'hC658, 16'hDF1A, 16'hCED9, 16'hD6DA, 16'hDF1A, 16'hB594, 16'hB513, 16'h9C50, 16'h7ACB, 16'hA450, 16'hD596, 16'hD596, 16'hC515, 16'hAC92, 16'hA451, 16'hA451, 16'h9C11, 16'hC5D7, 16'hDEDA, 16'hF79E, 16'hFFDF, 16'hEF5D, 16'h9CD2, 16'hAD54, 16'hD69A, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h9492, 16'h8C51, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'hA514, 16'h8C51, 16'h8C51, 16'h8C51, 16'hB596, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'hC618, 16'hDEDB, 16'hCE59, 16'h8C51, 16'h7B8E, 16'h9450, 16'hAD14, 16'hC596, 16'hCE17, 16'hD618, 16'hDE9A, 16'hBDD5, 16'h9D12, 16'hDF1B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hC618, 16'h9492, 16'h8410, 16'hF7DE, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h738E, 16'h634B, 16'h73CD, 16'h634B, 16'h5289, 16'h62CA, 16'h7B8D, 16'h8C50, 16'hB5D5, 16'hB5D6, 16'hB5D5, 16'hBE57, 16'hCE99, 16'hD6DA, 16'hDF1B, 16'hCE98, 16'hCE99,
        16'hCE99, 16'hAD95, 16'h5A89, 16'h1800, 16'h3000, 16'h000, 16'h000, 16'h000, 16'h041, 16'h2104, 16'h1082, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h1882, 16'h000, 16'h000, 16'h2104, 16'hC698, 16'hD75B, 16'hD71B, 16'hD75B, 16'hCF1A, 16'hBE16, 16'hC657, 16'hB594, 16'hAD13, 16'hA4D2, 16'h9450, 16'h9C91, 16'hA4D1, 16'h9450, 16'h8C0F, 16'h730B, 16'h8B8E, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h7BCF, 16'h8410, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hDEDB, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hD69A, 16'hB596, 16'hA513, 16'h840F, 16'h7BCE, 16'h840F, 16'h7BCE, 16'h6B8C, 16'h000, 16'h73CE, 16'hBE17, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD6DA, 16'hAD54, 16'h9C92, 16'h7BCE, 16'h7C0F, 16'hA595, 16'hBE57, 16'hC698, 16'hD6DA, 16'hDF5B, 16'hD6DA, 16'hC698, 16'hDF1B, 16'hD71B, 16'hD71B, 16'hD71A, 16'hD71A, 16'hD71B, 16'hB616, 16'hBE57, 16'hDF5B, 16'hDF9C, 16'hA554, 16'h000, 16'h1104, 16'h1083, 16'h2104, 16'h18C3, 16'h800, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h1041, 16'h1882, 16'h000, 16'h000, 16'h1881, 16'h734C, 16'h4A08, 16'hCE98, 16'hD71A, 16'hD71A, 16'hD71A, 16'hCED9, 16'hB615, 16'hD71A, 16'hDF1B, 16'hE71B, 16'hDF1A, 16'hE71B, 16'hE71B, 16'hDF1A, 16'hDF1A, 16'hE71B, 16'hDE99, 16'hC617, 16'h8C0F,
        16'h734C, 16'hB555, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hEF5D, 16'hE71C, 16'hE71C, 16'hDEDB, 16'hDEDB, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hBD96, 16'h738D, 16'h6B8D, 16'h9D12, 16'hB5D5, 16'hCED9, 16'hD71A, 16'hD71A, 16'hCF1A, 16'hCF1A,
        16'hCEDA, 16'hD71A, 16'hADD5, 16'hBE98, 16'hD71A, 16'hCEDA, 16'hCEDA, 16'hCEDA, 16'hCEDA, 16'hD71A, 16'hBE57, 16'hC698, 16'hD71A, 16'hD71A, 16'hAD95, 16'h000, 16'h18C3, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h1082, 16'h18C2, 16'h841, 16'h000, 16'h000, 16'h800, 16'h7B4D, 16'hCD95, 16'hC555, 16'h5289, 16'hD6D9, 16'hCEDA, 16'hCF1A, 16'hD71A, 16'hCE99, 16'hB616, 16'hCF1A, 16'hCEDA, 16'hD6DA, 16'hD6DA, 16'hD6D9, 16'hD71A, 16'hB616, 16'hC698, 16'hD71A, 16'hD71A, 16'hDF1B, 16'hDF1B, 16'hCE58, 16'h9C91, 16'h5A49, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h5289, 16'h73CD, 16'hB616, 16'hCED9, 16'hD71A, 16'hAE16, 16'hBE98, 16'hCED9, 16'hC6D9, 16'hCED9, 16'hC6D9, 16'hCEDA, 16'hC6D9, 16'h9D53, 16'hCED9, 16'hCEDA, 16'hCEDA, 16'hCEDA, 16'hCEDA, 16'hCEDA, 16'hD71A, 16'hADD6, 16'hBE57, 16'hD71B, 16'hDF5B, 16'hC658, 16'h000, 16'h18C2, 16'h18C2, 16'h1082, 16'h1041, 16'h1041, 16'h1041, 16'h1081, 16'h1082, 16'h1882, 16'h1882, 16'h1041, 16'h000, 16'h000, 16'h000, 16'h000, 16'h5208, 16'h93CF, 16'hC555, 16'hDE18, 16'hE659, 16'hBCD3, 16'h2984, 16'hCED9, 16'hDF5B, 16'hCEDA, 16'hD71A, 16'hCE98, 16'hB616,
        16'hCF1A, 16'hCEDA, 16'hCEDA, 16'hD6DA, 16'hD6D9, 16'hCED9, 16'hA554, 16'hCED9, 16'hD71A, 16'hD6DA, 16'hD6DA, 16'hD71A, 16'hDF1A, 16'hD6D9, 16'hCE59, 16'h840F, 16'h6B4D, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE99,
        16'h2983, 16'hAD95, 16'hD6DA, 16'hCED9, 16'hC699, 16'hCED9, 16'hAE16, 16'hA5D5, 16'hCF1A, 16'hCED9, 16'hC6D9, 16'hCED9, 16'hCEDA, 16'hC698, 16'hA594, 16'hCED9, 16'hCEDA, 16'hCEDA, 16'hCEDA, 16'hCEDA, 16'hCEDA, 16'hD71A, 16'hBE57, 16'hC698, 16'hCED9, 16'hB5D6, 16'h8450, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h000, 16'h2103, 16'h62CB, 16'h9410, 16'hBD54, 16'hD5D7, 16'hDE18, 16'hDE18, 16'hDE17, 16'hDE18, 16'hBD14, 16'h18C1, 16'h634C, 16'hADD5, 16'hD71B, 16'hD71B, 16'hCED9, 16'hB616, 16'hCF1A, 16'hCED9, 16'hCEDA, 16'hCED9, 16'hD71A, 16'hC657, 16'hAD95, 16'hD71A, 16'hD6D9, 16'hDF1A, 16'hDEDA, 16'hBDD6, 16'h9490, 16'h9CD2, 16'hB5D6, 16'hD699, 16'hA513, 16'h5A89, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h4207, 16'hADD6, 16'hD71A, 16'hC698, 16'hC698, 16'hC699, 16'hCED9, 16'hB617, 16'h9D95, 16'hCF1A, 16'hC6D9, 16'hC6D9, 16'hC6D9, 16'hCEDA, 16'hC699, 16'hA595, 16'hCEDA, 16'hCEDA, 16'hCEDA, 16'hCEDA, 16'hC6DA, 16'hD71B, 16'hC698, 16'h7C4F, 16'h5B4B, 16'h4288, 16'h5B0B, 16'h8C90, 16'h5289, 16'h838E, 16'h7B8D, 16'h62CA, 16'h5A89, 16'h5249, 16'h5A89, 16'h628A, 16'h730C, 16'h838E, 16'h9C51, 16'hBD14, 16'hCD95, 16'hDE17, 16'hDE18, 16'hDE18, 16'hDE17,
        16'hDE17, 16'hDE17, 16'hDE17, 16'hDE58, 16'hBD13, 16'h52C9, 16'hA552, 16'h4247, 16'h6BCE, 16'hC698, 16'hD6DA, 16'hBE57, 16'hCEDA, 16'hCED9, 16'hCEDA, 16'hCED9, 16'hD71A, 16'hB616, 16'hB616, 16'hD71A, 16'hDF1B, 16'hCE58, 16'h6B4C, 16'h5A89, 16'h6ACB, 16'h734C, 16'hC657, 16'hC698, 16'hDF1B, 16'h8C51, 16'h9C92, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h740F, 16'hD6DA, 16'hC6D9, 16'hCEDA, 16'hC699, 16'hC698, 16'hCED9, 16'hB617, 16'h9D94, 16'hCEDA, 16'hC6D9, 16'hC6D9, 16'hC6D9, 16'hCED9, 16'hC698, 16'h9D95, 16'hCED9, 16'hCEDA, 16'hCED9, 16'hC6D9, 16'hD71B, 16'hB616, 16'h52C9, 16'h9D12, 16'hAD95, 16'hC658, 16'hD6DA, 16'hDF1A, 16'h6B4C, 16'hCD95, 16'hE658, 16'hDE17, 16'hDE17, 16'hDDD7, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE18, 16'hE618, 16'hDE18, 16'hDE18, 16'hDE17, 16'hD5D7, 16'hD617, 16'hD617, 16'hD617, 16'hD617, 16'hD617, 16'hDE58, 16'hBD13, 16'h4A48, 16'hCE99, 16'hC698, 16'h7C0F, 16'h2103, 16'h94D2, 16'hC698, 16'hCEDA, 16'hCED9, 16'hCED9, 16'hCED9, 16'hD71A, 16'hA594, 16'hBE57, 16'hE75B, 16'hB595, 16'h3945, 16'h9450, 16'hD658, 16'hD69A, 16'hA514, 16'h9D13, 16'hD6DA, 16'hD699, 16'hCE99, 16'h5ACA, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h738D, 16'hB5D6, 16'hCEDA, 16'hB5D6, 16'hA594, 16'hC699, 16'hC699, 16'hCED9, 16'hB657, 16'h9D54, 16'hCED9, 16'hC6D9, 16'hC6D9, 16'hC6D9, 16'hCED9, 16'hC698, 16'h9D94, 16'hCED9, 16'hCEDA, 16'hC6D9, 16'hD71A, 16'hADD6, 16'h31C6, 16'hB5D5, 16'hCE98, 16'hC617, 16'hB5D5, 16'h9491, 16'h8C50, 16'h39C6, 16'hBD14, 16'hE618, 16'hDE17, 16'hDE18,
        16'hDE18, 16'hDE18, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hD617, 16'hD617, 16'hD617, 16'hDE18, 16'hC514, 16'h39C6, 16'hA594, 16'hC699, 16'hCEDA, 16'hAD94, 16'h000, 16'h8C91, 16'hD71A, 16'hCED9, 16'hCED9, 16'hCEDA, 16'hCED9, 16'h9D53, 16'hD6DA, 16'hA553, 16'h41C5, 16'hBD95, 16'hDEDA, 16'hD699, 16'hCE99, 16'hD6DA, 16'h8C91, 16'hB5D6, 16'hD6DA, 16'hDF1A, 16'h840F, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hA514, 16'hA514, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h630C, 16'hCE99, 16'hADD6, 16'h8C91, 16'h7C0F, 16'h6B8D, 16'hC698, 16'hCED9, 16'hBE58, 16'h9594, 16'hCED9, 16'hC6D9, 16'hC6D9, 16'hC6D9, 16'hCED9, 16'hC6D9, 16'hA595, 16'hC6D9, 16'hC6D9, 16'hD71A, 16'hB616, 16'h1942, 16'hAD95, 16'hD6DA, 16'h8C50, 16'h000, 16'h31C5, 16'h39C5, 16'h4A47, 16'h3144, 16'hC555, 16'hDE18, 16'hDE17, 16'hDE18, 16'hDE18, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hD617, 16'hDE18, 16'hC554, 16'h20C2, 16'h4A88, 16'h8450, 16'hBE17, 16'hBE16, 16'hB5D5, 16'h1000, 16'h9D54, 16'hD71A, 16'hCED9, 16'hCF1A, 16'hC698, 16'hAD95, 16'h9D13, 16'h39C6, 16'hC617, 16'hDE9A, 16'hCE99, 16'hD699, 16'hCE99, 16'hD6DA, 16'hC658, 16'h8C91, 16'hD6D9, 16'hDF1B, 16'hA513, 16'hAD54,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8410, 16'h8410, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h6B8D, 16'hCE99, 16'h8C91, 16'hCE99, 16'hDEDA, 16'h9491, 16'h6B8D, 16'hCEDA, 16'hBE58, 16'h9553, 16'hC6D9, 16'hC6D9, 16'hC6D9, 16'hC6D9, 16'hCED9, 16'hC6D9, 16'h9D94, 16'hC699, 16'hD71B, 16'hAE16, 16'h3A06, 16'hB595,
        16'hD699, 16'hD699, 16'h9CD2, 16'h31C4, 16'h630A, 16'h5ACA, 16'h4A48, 16'h3986, 16'hCD96, 16'hDE18, 16'hDE17, 16'hDE18, 16'hDE18, 16'hDE18, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE18, 16'hC554, 16'h2903, 16'h5AC9, 16'h4A88, 16'h7BCD, 16'h740D, 16'hCE58, 16'hB595, 16'h000, 16'hB616, 16'hD71A, 16'hCF1A, 16'hC698, 16'h634C, 16'h6B4C, 16'hCE58, 16'hD69A, 16'hD699, 16'hD699, 16'hD699, 16'hD699, 16'hCE99, 16'hD6DA, 16'h94D2, 16'hC617, 16'hE71B, 16'hB595, 16'h9491, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8C51, 16'h8C51, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBE17, 16'h8C91, 16'hB5D6, 16'hA554, 16'hDEDA, 16'hD699, 16'hDF1A, 16'h8450, 16'h9513, 16'hCEDA, 16'h9513, 16'hC6D9, 16'hC6D9, 16'hC6D9, 16'hC6D9, 16'hC6D9, 16'hCED9, 16'h9554, 16'hCEDA, 16'hB616, 16'h000, 16'hAD54, 16'hD699, 16'hC658, 16'hD699, 16'hB595, 16'h39C6, 16'h4A48, 16'h41C6, 16'h2800, 16'h8B8E, 16'hDE18, 16'hDDD7, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hCD95, 16'h3144, 16'h5AC9, 16'h4206, 16'h5ACA, 16'hC616, 16'hCE58, 16'hD699, 16'h9491, 16'h000, 16'hBE57, 16'hD6D9, 16'h73CE, 16'h6B4C, 16'hD658, 16'hD699,
        16'hCE99, 16'hD699, 16'hD699, 16'hD699, 16'hD699, 16'hCE99, 16'hD6DA, 16'hAD95, 16'hAD95, 16'hE71B, 16'hBDD6, 16'h840F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h9D13, 16'h9D13, 16'hC617, 16'hD6D9, 16'hD699, 16'hD6D9, 16'hCE99, 16'h4A49, 16'hB617, 16'hA594,
        16'hBE98, 16'hC6D9, 16'hC6D9, 16'hC6D9, 16'hC6D9, 16'hCED9, 16'hA5D6, 16'hA594, 16'h2985, 16'hA553, 16'hCE99, 16'hCE58, 16'hCE58, 16'hD699, 16'hC617, 16'h3185, 16'h5A48, 16'h93CE, 16'h7B0B, 16'hCD95, 16'hDE18, 16'hDDD7, 16'hDDD7, 16'hDDD7, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hD5D7, 16'hDE17, 16'hDDD7, 16'h5208, 16'h000, 16'h6B4C, 16'hC617, 16'hD698, 16'hCE58, 16'hCE58, 16'hCE98, 16'h7BCE, 16'h5289, 16'h5ACB, 16'h6B0B, 16'hCE17, 16'hDE99, 16'hCE99, 16'hCE99, 16'hD699, 16'hD699, 16'hCE99, 16'hCE99, 16'hCE99, 16'hD6DA, 16'hBE17, 16'h94D2, 16'hDF1B, 16'hC658, 16'h73CE, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h9492, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h8C51, 16'h94D2, 16'h9D13, 16'hCE99, 16'hD699, 16'hD699, 16'hCE58, 16'hD6DA, 16'hAD95, 16'h630C, 16'hA594, 16'hBE57, 16'hCED9, 16'hC6D9, 16'hC6D9, 16'hC6D9, 16'hD75B, 16'h9513, 16'h000, 16'hAD94, 16'hD699, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hD658, 16'h6B4C, 16'hA450, 16'hAC51, 16'hC554, 16'hDE18, 16'hDDD7, 16'hDDD7, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hD617, 16'hD5D7, 16'hDE18, 16'hDE18, 16'hA491, 16'h20C1, 16'h8C50, 16'hCE58,
        16'hD698, 16'hCE58, 16'hD658, 16'hCE98, 16'hDED9, 16'hC617, 16'h000, 16'h6B0C, 16'hAD14, 16'hAD13, 16'hAD13, 16'hD699, 16'hD699, 16'hCE99, 16'hCE99, 16'hCE99, 16'hCE99, 16'hCE99, 16'hD6DA, 16'hC658, 16'h94D2, 16'hD6DA, 16'hCE99, 16'h6B4C, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hEF5D, 16'hE71C, 16'hE71C, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hE71C, 16'h9CD3, 16'h9492, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'h8410, 16'h8C50, 16'hA554, 16'hD699, 16'hEF1C, 16'hFF5E, 16'hEF1D, 16'hD699, 16'hD6D9, 16'h7C0F, 16'h530A, 16'hC658, 16'hCEDA, 16'hC6D9, 16'hCED9, 16'hCF1A, 16'hA594, 16'h000, 16'h8C50, 16'hD699, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hD699, 16'h9492, 16'h834C, 16'hCD96, 16'hDDD7, 16'hDDD7, 16'hDDD7, 16'hDDD7, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hD617, 16'hD617, 16'hDE17, 16'hDE17, 16'hDE17, 16'hD617, 16'hD5D7, 16'hDE17, 16'hDE58, 16'hC554, 16'h628A, 16'h62CB, 16'hBDD5, 16'hD699, 16'hCE98, 16'hCE58, 16'hCE58, 16'hD698, 16'hDE99, 16'hAD54, 16'h3986, 16'hA513, 16'hD699, 16'hD699, 16'hDEDA, 16'hBDD6, 16'hAD54, 16'hD6DA, 16'hCE99, 16'hCE99, 16'hCE99, 16'hCED9, 16'hCE99, 16'hD6D9, 16'hCE99, 16'h94D2, 16'hCE99, 16'hD6DA, 16'h6B8D, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'hAD55, 16'h8C51, 16'h8C51, 16'h8C51, 16'h8C51, 16'hB596, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hB596, 16'h9492, 16'h8C51, 16'h9492, 16'h9492, 16'h8410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h7BCF, 16'h840F, 16'hBDD6, 16'hD699, 16'hF75E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hBD55, 16'hB554, 16'h6B0C, 16'h7C0F, 16'hD71A, 16'hCED9, 16'hCF1A, 16'h8CD2, 16'h4A08, 16'h8C50, 16'h9491, 16'hD699, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hD699, 16'hC617, 16'h6289, 16'hCD96, 16'hDDD7, 16'hD5D7, 16'hDDD7, 16'hDDD7, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hD617, 16'hD617, 16'hD617, 16'hD617,
        16'hDE17, 16'hD5D7, 16'hD617, 16'hDE18, 16'hCDD6, 16'h8BCE, 16'h4207, 16'h9CD2, 16'hD658, 16'hD699, 16'hCE58, 16'hCE58, 16'hCE98, 16'hD699, 16'hD698, 16'h7BCE, 16'h5ACA, 16'hC5D6, 16'hDEDA, 16'hD699, 16'hD699, 16'hD699, 16'hD6DA, 16'h9CD2, 16'hC658, 16'hD69A, 16'hCE99, 16'hCED9, 16'hCE99, 16'hCE99, 16'hCED9, 16'hD6DA, 16'h94D2, 16'hC658, 16'hD6DA, 16'h738E, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hAD55, 16'h8410, 16'h8C51, 16'h9492, 16'h8C51, 16'h9492, 16'h9492, 16'h8410, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hDEDB, 16'hD69A, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8410, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'h9492, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF9D, 16'h5B0B, 16'h840F, 16'hC617, 16'hD699, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hDE9B, 16'hC5D7, 16'hFFDF, 16'hEF1C, 16'h62CB, 16'h8C91, 16'hCED9, 16'h740E, 16'h3185, 16'hC617, 16'hAD54, 16'h840F, 16'hD699, 16'hCE58, 16'hCE58, 16'hCE59, 16'hCE59, 16'hCE59, 16'hCE58, 16'hD699, 16'h7BCE, 16'hAC51, 16'hDE18, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD617, 16'hDE17, 16'hDE17, 16'hDE17, 16'hDE17, 16'hD617, 16'hD617, 16'hD617, 16'hD5D7, 16'hD5D7, 16'hDE18, 16'hD617, 16'hA451, 16'h4A07, 16'h8C50, 16'hCE17, 16'hD699, 16'hD658, 16'hCE58, 16'hCE58, 16'hD698, 16'hDE99, 16'hB595, 16'h5249, 16'h9451, 16'hD699, 16'hDEDA, 16'hD699, 16'hD699, 16'hD699, 16'hD699, 16'hDEDA, 16'hB595, 16'hAD54, 16'hD6DA, 16'hCE99, 16'hCED9, 16'hCE99, 16'hCE99, 16'hCED9, 16'hD6DA, 16'h9D13, 16'hB616, 16'hDF1B, 16'h7C0F, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9CD3, 16'h8410, 16'h9492, 16'h9492, 16'h8C51, 16'hA514, 16'hA514, 16'h8C51, 16'h9492, 16'h8410, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hBDD7, 16'h9492, 16'h8C51, 16'h8410, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h9492, 16'h9492, 16'h8410, 16'h9CD3, 16'h9CD3, 16'h9492,
        16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h4207, 16'h94D2, 16'hCE58, 16'hD699, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hB555, 16'hF75D, 16'hFF9F, 16'hFF9F, 16'hF75D, 16'h8C10, 16'h000, 16'h5ACA, 16'hBDD6, 16'hCE58, 16'hB595, 16'h73CE, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE98, 16'hCE58, 16'hD699, 16'hBDD6, 16'h5A07, 16'hD596, 16'hDE17,
        16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD617, 16'hD617, 16'hD617, 16'hD617, 16'hD617, 16'hD617, 16'hD5D7, 16'hD5D7, 16'hDE17, 16'hDE17, 16'hB4D3, 16'h6289, 16'h630C, 16'hBDD6, 16'hDE99, 16'hD658, 16'hCE58, 16'hCE58, 16'hD698, 16'hDED9, 16'hCE57, 16'h738D, 16'h5ACA, 16'hBD96, 16'hDEDA, 16'hD699, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE98, 16'hD6D9, 16'hCE58, 16'h9491, 16'hD699, 16'hCE99, 16'hCE99, 16'hCE99, 16'hD699, 16'hCE99, 16'hD6DA, 16'hA554, 16'hB5D6, 16'hD71A, 16'hAD95, 16'h8C50, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h7BCF, 16'h9CD3, 16'h9492, 16'h8C51, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8C51, 16'h9492, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h9CD3, 16'h8410, 16'h9492, 16'h9492, 16'h9CD3, 16'h8410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h9492, 16'h8C51, 16'hA514, 16'hDEDB, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h9CD3, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE58, 16'h1080, 16'hAD54, 16'hCE99, 16'hD69A, 16'hFF9F, 16'hFFDF, 16'hE6DB, 16'hC5D7, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9E, 16'h8C10, 16'h6B4C, 16'hC5D6, 16'hCE58, 16'hC617, 16'h738D, 16'hC658, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE98, 16'hCE98, 16'hCE98, 16'hD699, 16'h83CF, 16'h7289, 16'hDDD7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD617, 16'hD5D7, 16'hD617, 16'hD5D7, 16'hD5D7, 16'hDE17, 16'hC554, 16'h72CA, 16'h5ACA, 16'hAD54, 16'hD699, 16'hD699, 16'hCE58, 16'hCE58, 16'hD698, 16'hD6D9, 16'hCE58, 16'h8C50, 16'h5289, 16'hA4D2, 16'hCE18, 16'hD658, 16'hD699, 16'hCE58, 16'hD659, 16'hE6DB, 16'hF75D, 16'hF75D, 16'hDEDA, 16'hCE98, 16'hD6D9, 16'h9C92, 16'hC658, 16'hD699, 16'hCE99, 16'hCE99, 16'hD699, 16'hCE99, 16'hD6DA,
        16'hADD5, 16'hAD95, 16'hD6DA, 16'hC698, 16'h3A07, 16'h9CD3, 16'hDEDB, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9CD3, 16'h8C51, 16'h9492, 16'h8410, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h8C51, 16'h9492, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'hBDD7,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hD69A, 16'hEF5D, 16'hFFDF, 16'hF79E, 16'hA514, 16'h8410, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hA514, 16'h4A49, 16'h4A49, 16'hC617, 16'hCE58, 16'hDE9A, 16'hFF9F, 16'hFFDF, 16'hBD96, 16'hE6DB, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'h9492, 16'h18C0, 16'hB595, 16'hD699, 16'h738D,
        16'hBDD6, 16'hD699, 16'hCE58, 16'hCE58, 16'hCE59, 16'hCE99, 16'hCE99, 16'hCE99, 16'hD699, 16'hCE58, 16'h4A08, 16'h8B8D, 16'hE617, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hD5D7, 16'hDE18, 16'hCDD6, 16'h838D, 16'h5A8A, 16'h9CD2, 16'hCE58, 16'hD699, 16'hCE58, 16'hCE58, 16'hD699, 16'hDED9, 16'hCE58, 16'h9CD2, 16'h5ACA, 16'h840F, 16'hCE18, 16'hE6DA, 16'hEEDB, 16'hAD13, 16'hD659, 16'hF75D, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hDEDA, 16'hD699, 16'hA513, 16'hB596, 16'hD6DA, 16'hCE99, 16'hD699, 16'hD699, 16'hCE99, 16'hD6D9, 16'hBE17, 16'hA594, 16'hCED9, 16'hCED9, 16'h9512, 16'h4207, 16'h4A48, 16'h4208, 16'h9492, 16'hC618, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB596, 16'h8C51, 16'h8410, 16'hCE59, 16'hFFDF, 16'hEF5D, 16'hA514, 16'h8C51, 16'h8C51, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8410, 16'h9492, 16'h8410, 16'hD69A, 16'hCE59, 16'h8C51, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8C51, 16'h8C51, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8C51, 16'h8C51, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hAD55, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h7BCF, 16'h9492, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9CD3, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'hCE59, 16'hA514, 16'h8410, 16'h3185, 16'h630B, 16'h2945, 16'h840F, 16'hD699, 16'hCE58, 16'hDE9A, 16'hFF9F, 16'hFF5E, 16'hB555, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hF75D, 16'hAD14, 16'h4207, 16'hB595, 16'h9491, 16'hA513, 16'hD699, 16'hCE58, 16'hCE58, 16'hCE59, 16'hCE99, 16'hCE99, 16'hCE99, 16'hCE58, 16'hD699, 16'hC617, 16'h5A89, 16'h9BCE, 16'hD5D6, 16'hDDD7, 16'hD5D7, 16'hDDD7, 16'hDE18, 16'hDE18, 16'hD5D7, 16'hA491, 16'h6289, 16'h9451, 16'hCE58, 16'hD699, 16'hCE58, 16'hCE58, 16'hD699, 16'hD699, 16'hCE58, 16'h9451, 16'h41C6, 16'h734D, 16'hCE17, 16'hE6DB, 16'hEF1C, 16'hF75D, 16'hFFDF, 16'hD618, 16'hD619, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFFDF, 16'hEF1C, 16'hD699, 16'hB595, 16'hAD54, 16'hD6DA, 16'hCE99, 16'hD699, 16'hD699, 16'hCE99, 16'hCE99, 16'hBE17, 16'hA553, 16'hCE99, 16'hC698, 16'hC658, 16'hA553, 16'h7BCE, 16'h630B, 16'h8C50, 16'h634B, 16'h4A48, 16'h738D, 16'hB595, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8410, 16'h9492, 16'hA514, 16'hAD55, 16'h8C51, 16'h8C51, 16'h9492, 16'h8410, 16'hDEDB, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h9492, 16'h8C51, 16'hC618, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h9CD3, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8C51, 16'h8C51, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8C51, 16'h8C51, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9CD3, 16'h8410, 16'h8410, 16'hF79E, 16'hEF5D, 16'h8410, 16'h9CD3, 16'h8410, 16'hE71C, 16'hEF5D, 16'h7BCF, 16'h8C51, 16'h8410, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hC618, 16'h840F, 16'h630B, 16'h630B, 16'h840F, 16'h8C50, 16'h8C51, 16'hAD14, 16'h000, 16'hAD54, 16'hD699, 16'hCE58, 16'hD699, 16'hFFDF, 16'hE69B, 16'hC596,
        16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF5E, 16'h8BCF, 16'h3185, 16'h4A88, 16'h9CD2, 16'hDEDA, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE59, 16'hCE59, 16'hCE58, 16'hCE98, 16'hD699, 16'hCE58, 16'h83CE, 16'h000, 16'h8B8D, 16'hDDD7, 16'hDE17, 16'hD5D7, 16'hC555, 16'hBD14, 16'h8BCF, 16'h83CF, 16'hBDD6, 16'hD699, 16'hD658, 16'hD658, 16'hD699, 16'hD699, 16'hC5D6, 16'h840F, 16'h5207, 16'h8C0F, 16'hD659, 16'hF75E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hEF1D, 16'hBD55, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF75D, 16'hD699, 16'hC617, 16'h9CD2, 16'hD699, 16'hD699, 16'hD699, 16'hCE99, 16'hCE59, 16'hCE99, 16'hC658, 16'hA553, 16'hC698, 16'hC658, 16'hC657, 16'hC658, 16'hA553, 16'h39C6, 16'hBE17, 16'hD6DA, 16'hC617, 16'hA554, 16'h7BCE, 16'h3185, 16'h5B0B, 16'hAD55, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8410, 16'h9492, 16'h8C51, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'h9CD3, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h9492, 16'hF79E, 16'hFFDF, 16'hEF5D, 16'h9492, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8C51, 16'h8C51, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9CD3, 16'h9492, 16'h8C51, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9CD3, 16'h8410, 16'hDEDB, 16'hFFDF, 16'h9492, 16'h7BCF, 16'h9CD3, 16'hF79E, 16'hFFDF, 16'hD69A, 16'hB596, 16'hE71C,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'hAD55, 16'h528A, 16'h18C1, 16'h8C51, 16'hA513, 16'hA4D3, 16'hAD14, 16'hBDD6, 16'hA4D2, 16'h000, 16'h5ACA, 16'hBDD6, 16'hD699, 16'hD658, 16'hD659, 16'hFF9F, 16'hCDD8, 16'hD659, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE9A, 16'hCDD8, 16'hDE9A, 16'h6B0C, 16'h3185, 16'hAD54, 16'hD699, 16'hD699, 16'hD699, 16'hCE59, 16'hCE58, 16'hD699, 16'hD699, 16'h9CD2, 16'h4207, 16'h7BCF, 16'hC617, 16'h630B, 16'h9C0F, 16'hE658, 16'h730C, 16'h5A8A, 16'h4A08, 16'h49C6, 16'hC5D7, 16'hDE9A, 16'hD699, 16'hD699, 16'hCE17, 16'h9CD2, 16'h5A89, 16'h5208, 16'hA4D3, 16'hE6DB, 16'hFFDF, 16'hFFDF,
        16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hB514, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hDE99, 16'hCE58, 16'h9491, 16'hD699, 16'hD699, 16'hD699, 16'hCE58, 16'hCE59, 16'hCE58, 16'hCE58, 16'hA553, 16'hBE17, 16'hC657, 16'hC657, 16'hCE98, 16'h7BCE, 16'h52C9, 16'h9D12, 16'hA513, 16'hBDD6, 16'hCE99, 16'hD699, 16'hCE58, 16'hA513, 16'h4A89, 16'h000, 16'h7BCF, 16'hBDD6, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hEF5D, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'h8410, 16'h8410, 16'h8410, 16'h9492, 16'h8C51, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hD69A, 16'h8C51, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8C51, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h8C51, 16'hC618, 16'hF79E, 16'hDEDB, 16'h9CD3, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA514, 16'h7BCF, 16'hA514, 16'hF79E, 16'hFFDF, 16'hE71C, 16'hC618, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h840F, 16'h5289, 16'h9491, 16'h738D, 16'h9CD2, 16'hBD95, 16'hB595, 16'hC617,
        16'hD659, 16'hD699, 16'hCE18, 16'h2104, 16'h9C91, 16'hCE58, 16'hD659, 16'hD658, 16'hD659, 16'hFF5E, 16'hBD56, 16'hE6DC, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hBD96, 16'hFF9E, 16'hFFDF, 16'hF71D, 16'hB555, 16'h62CB, 16'h630B, 16'h9CD2, 16'hC617, 16'hCE58, 16'hD699, 16'hCE58, 16'h7BCE, 16'h630C, 16'hB595, 16'hCE58, 16'hCE58, 16'hB595, 16'h5248, 16'h940F, 16'h4A07, 16'hCE18, 16'hCE17, 16'h8C0F, 16'h5249, 16'hBD95, 16'hA4D2, 16'h7B8D, 16'h5A89, 16'h730C, 16'hC596, 16'hDE59, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hBD56, 16'hE6DB, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hE6DB, 16'hCE58, 16'h9CD2, 16'hCE58, 16'hD699, 16'hCE59, 16'hCE58, 16'hCE58, 16'hCE58, 16'hD699, 16'hAD54, 16'hB5D6, 16'hC658, 16'hC658, 16'h7BCE, 16'h738E, 16'hC617, 16'hC617, 16'hA513, 16'h9491, 16'h8C90, 16'hB5D6, 16'hD699, 16'hD699, 16'hD699, 16'h7BCE, 16'h9CD2, 16'h8C50, 16'h5ACA,
        16'h8C51, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9CD3, 16'h9492, 16'h8C51, 16'hBDD7, 16'hDEDB, 16'hE71C, 16'hC618, 16'h9492, 16'h9492, 16'h8410, 16'hBDD7, 16'hFFDF, 16'hD69A, 16'h8C51, 16'h8C51, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8410, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8410, 16'h9CD3, 16'h8C51, 16'h8C51, 16'h8410, 16'h9492, 16'h9492, 16'h8410, 16'h8C51, 16'h7BCF, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E,
        16'hDEDB, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDE, 16'hC618, 16'h6B4C, 16'h630B, 16'hA513, 16'hD658, 16'hE6DA, 16'h7B8D, 16'hA513, 16'hD699, 16'hD699, 16'hD659, 16'hD699, 16'hD699, 16'hD699, 16'h6B0B, 16'hB554, 16'hDE9A, 16'hD658, 16'hD659, 16'hD659, 16'hF71D, 16'hB514, 16'hF71D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE6DB, 16'hCDD8, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9E, 16'hE6DC, 16'hBD96, 16'h7BCE, 16'h62CB, 16'h528A, 16'h738D, 16'h2102, 16'h5ACA, 16'hC617, 16'hC617, 16'hC617, 16'hCE57, 16'hD658, 16'h738D, 16'h000, 16'h9C51, 16'hB554, 16'h8C0F, 16'h5A49,
        16'h4186, 16'h730C, 16'hA493, 16'hCDD8, 16'hEF1D, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'hD659, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD619, 16'hD618, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE71C, 16'hD699, 16'h9C92, 16'hC617, 16'hD699, 16'hCE58, 16'hCE58, 16'hD658, 16'hD658, 16'hD699, 16'hBDD6, 16'hAD54, 16'hD699, 16'h738D, 16'h738D, 16'hCE59, 16'hCE58, 16'hCE58, 16'hD659, 16'hCE58, 16'hBDD7, 16'h9491, 16'hAD54, 16'hD699, 16'hC617, 16'h73CD, 16'hCE58, 16'hDEDA, 16'hCE58, 16'h9CD2, 16'h5ACA, 16'h734D, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD55, 16'h8C51, 16'h8410, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8C51, 16'h8C51, 16'hAD55, 16'hFFDF, 16'hDEDB, 16'h8C51, 16'h9492, 16'h9492, 16'hE71C, 16'hFFDF, 16'hF79E, 16'hA514, 16'h8C51, 16'h9492, 16'h8410, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hA514, 16'h8410, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'h8C51, 16'hCE59, 16'hC618, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7,
        16'h630B, 16'h6B4C, 16'hBD95, 16'hD659, 16'hDE9A, 16'hD659, 16'hD699, 16'h840F, 16'hA4D2, 16'hDE99, 16'hCE58, 16'hD699, 16'hCE17, 16'hAD13, 16'hA513, 16'h630B, 16'h9C91, 16'hDE9A, 16'hD659, 16'hD699, 16'hD659, 16'hEEDB, 16'hB514, 16'hF75D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hCE18, 16'hDE9B, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hEF1C, 16'hBD55, 16'hAD14, 16'hA4D3, 16'h8C10, 16'h6B4C, 16'h6B0B, 16'h5289, 16'h6B0C, 16'h630B, 16'h3944, 16'h4A07, 16'h7B4D, 16'h83CF, 16'hA4D3, 16'hCE18, 16'hEF1C, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hD619, 16'hF71D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE6DB, 16'hBD96, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF75D, 16'hD699, 16'hA513, 16'hBDD6, 16'hD699, 16'hCE58, 16'hD658, 16'hD658, 16'hD658, 16'hCE58, 16'hCE18, 16'hB555, 16'h83CF, 16'h5ACA, 16'hCE58, 16'hD659, 16'hCE58,
        16'hCE58, 16'hCE58, 16'hCE58, 16'hD658, 16'hD699, 16'h9CD3, 16'hB5D5, 16'h840F, 16'hB555, 16'hD699, 16'hCE58, 16'hD699, 16'hDE9A, 16'hD699, 16'hB595, 16'h6B4C, 16'h528A, 16'hBDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBDD7, 16'h8C51, 16'h8C51, 16'hC618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h8C51, 16'h8C51, 16'hB596, 16'hFFDF, 16'hF79E, 16'h9492, 16'h9492, 16'h9492, 16'h9492, 16'hB596, 16'h9492, 16'h8C51, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hC618, 16'h9CD3,
        16'h9492, 16'h9492, 16'hB596, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h738E, 16'h62CA, 16'hBD95, 16'hDE99, 16'hDE99, 16'hD658, 16'hD658, 16'hD659, 16'hDE99, 16'hAD54, 16'h83CF, 16'hDE99, 16'hD699, 16'hB555, 16'h9451, 16'hB555, 16'hD659, 16'hB555, 16'h6B4C, 16'hDE99, 16'hD699, 16'hD659, 16'hD659, 16'hDE59, 16'hACD3, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hC597, 16'hF75D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'hE69A, 16'hFFDF, 16'hFFDF,
        16'hFF9E, 16'hF75D, 16'hEF1C, 16'hDE9A, 16'hDE9A, 16'hDE9A, 16'hE6DB, 16'hEF1D, 16'hE69B, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE69B, 16'hE69A, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1D, 16'hACD3, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hFF9E, 16'hF75D, 16'hDE99, 16'hAD14, 16'hB554, 16'hD699, 16'hD658, 16'hD658, 16'hD658, 16'hCE58, 16'hCE58, 16'hD659, 16'h83CF, 16'h62CB, 16'hAD14, 16'h8C50, 16'hAD54, 16'hD699, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hD699, 16'h9491, 16'h9491, 16'hDE9A, 16'hD659, 16'hD699, 16'hD699, 16'hD659, 16'hD699, 16'hD699, 16'hDE99, 16'hBD96, 16'h5289, 16'h5ACB, 16'hD699, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h8410, 16'h8C51, 16'hB596, 16'hFFDF, 16'hF79E, 16'hCE59, 16'h8C51, 16'h9492, 16'h8410, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hCE59, 16'h7BCF, 16'h9492, 16'h9492, 16'h8C51, 16'h9492, 16'h9492, 16'h8C51, 16'h9492, 16'h8410, 16'h8C51, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD96, 16'h3903, 16'hAD13, 16'hDE99, 16'hDE99, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hD699, 16'hC617, 16'h630B, 16'hCE18, 16'hAD13, 16'hA513, 16'hD658, 16'hDE99, 16'hD659, 16'hD658, 16'h62CB, 16'hC5D7, 16'hDE99, 16'hD658, 16'hD659, 16'hCDD7, 16'hACD3, 16'hFF5E, 16'hF75E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hBD56, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'hDE9A, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD618, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF71D, 16'hD619, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hACD3, 16'hFF5E, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hEF1C, 16'hDE99, 16'hBD96, 16'hA4D2, 16'hD699,
        16'hD658, 16'hD658, 16'hCE58, 16'hD658, 16'hD658, 16'h7B8E, 16'h840F, 16'hD659, 16'hD659, 16'hC617, 16'h9C92, 16'h9491, 16'hCE58, 16'hD659, 16'hCE58, 16'hCE58, 16'hD699, 16'hBDD6, 16'h840F, 16'hD699, 16'hD699, 16'hD659, 16'hD699, 16'hD659, 16'hD699, 16'hD659, 16'hD658, 16'hD658, 16'hD699, 16'hD699, 16'hB555, 16'h5249, 16'h9451, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C51, 16'h9492, 16'h9CD3, 16'hB596, 16'h9CD3, 16'h8410, 16'h9492, 16'h8C51, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8C51, 16'h8C51, 16'h8C51,
        16'h8C51, 16'h9492, 16'hD69A, 16'hF79E, 16'hD69A, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h8C10, 16'h6ACA, 16'hDE59, 16'hEEDB, 16'hDE99, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hD699, 16'h7B8D, 16'h8C10, 16'hBDD6, 16'hD699, 16'hD658, 16'hD658, 16'hD658, 16'hDE99, 16'h83CF, 16'h9C91, 16'hDE9A, 16'hD659, 16'hDE99, 16'hBD55, 16'hACD3, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hEF1D, 16'hBD56,
        16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE6DB, 16'hE69B, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hD618, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'hCDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD14, 16'hEF1D, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hEF1C, 16'hDE59, 16'hCE17, 16'h9C92, 16'hD659, 16'hD658, 16'hD658, 16'hD659, 16'hC617, 16'h62CB, 16'h8C50, 16'hD699, 16'hD658, 16'hCE58, 16'hD659, 16'hD699, 16'hB555, 16'h8C10, 16'hC617, 16'hD659, 16'hCE58, 16'hC617, 16'h738D, 16'hC617, 16'hD699, 16'hD659, 16'hD699, 16'hD699, 16'hD699, 16'hD699, 16'hD659, 16'hD699, 16'hD699, 16'hCE58, 16'hCE58, 16'hD699, 16'hD658, 16'h8C50, 16'h31C6, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h9492, 16'h9492, 16'h9492, 16'h8C51, 16'h9492, 16'h9492, 16'h8410, 16'h9492, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'hDEDB, 16'hDEDB, 16'hE71C, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h83CE, 16'h940F, 16'hFF9E, 16'hFF9F, 16'hFF5D, 16'hFF9D, 16'hE6DB, 16'hDE99, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hD659, 16'hDE99, 16'hA513, 16'h738D, 16'hDE99, 16'hD658, 16'hD658, 16'hD658, 16'hD658, 16'hDE59, 16'hC5D6, 16'h734D, 16'hDE59, 16'hDE59, 16'hDE9A, 16'hB514, 16'hB514, 16'hFF5E, 16'hFF5D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFFDF, 16'hE6DB, 16'hC5D7, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE69B, 16'hEEDC, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD618, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hC597, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF,
        16'hBD56, 16'hE69A, 16'hFF9F, 16'hFF5D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hEEDB, 16'hDE59, 16'hD659, 16'h9C92, 16'hD618, 16'hD658, 16'hDE99, 16'hC5D6, 16'h5249, 16'hA4D3, 16'hDE99, 16'hD658, 16'hD658, 16'hD658, 16'hD658, 16'hCE58, 16'hD699, 16'hBDD6, 16'h9451, 16'hCE58, 16'hD699, 16'h83CF, 16'hB595, 16'hDE99, 16'hD659, 16'hD699, 16'hD699, 16'hD699, 16'hD699, 16'hD699, 16'hD659, 16'hD658, 16'hD658, 16'hCE58, 16'hCE58, 16'hD659, 16'hD699, 16'hE6DB, 16'hBDD6, 16'h4A08, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF79E, 16'h9492, 16'h8410, 16'h8C51, 16'h8C51, 16'h8C51,
        16'h9CD3, 16'hBDD7, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h8BCF, 16'hA492, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hF75D, 16'hDE9A, 16'hD658, 16'hD659, 16'hD659, 16'hD659, 16'hDE99, 16'hCE17, 16'h5A8A, 16'hCE17, 16'hD659, 16'hD658, 16'hD658, 16'hD618, 16'hDE99, 16'hCE17, 16'h41C7, 16'hBD96, 16'hDE9A,
        16'hE6DA, 16'hB514, 16'hBD15, 16'hF75D, 16'hFF5D, 16'hFF5D, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFFDF, 16'hD659, 16'hCE18, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE69A, 16'hEEDC, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hCE18, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hCDD7, 16'hF75D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hC5D7, 16'hD618, 16'hFF9E, 16'hFF5D, 16'hFF5E, 16'hFF5E, 16'hFF5D, 16'hDE5A, 16'hDE59, 16'hDE99, 16'hA492, 16'hC5D7, 16'hDE9A, 16'hB554, 16'h5248, 16'hBD96, 16'hDE9A, 16'hD658, 16'hD658, 16'hD658, 16'hCE58, 16'hCE58, 16'hD658, 16'hCE58, 16'hD699, 16'hBDD6, 16'hB595, 16'h9491, 16'h9CD2, 16'hDEDA, 16'hD658, 16'hD699, 16'hD659, 16'hD659, 16'hD699, 16'hD659, 16'hD658, 16'hD658, 16'hD699, 16'hDE99, 16'hE6DB, 16'hEEDC, 16'hF71D, 16'hF75D,
        16'hF75E, 16'hFFDF, 16'hE6DB, 16'h3903, 16'hCE58, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'hAD55, 16'hBDD7, 16'hCE59, 16'hE71C, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9451, 16'hA451, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hE6DB, 16'hD658, 16'hD659, 16'hD659, 16'hD659, 16'hDE99, 16'h738D, 16'hAD14, 16'hDE99, 16'hD658, 16'hD658, 16'hD659, 16'hACD3, 16'h838E, 16'h8C10, 16'h734D, 16'hDE99, 16'hE69A, 16'hB4D3, 16'hC556, 16'hEEDC, 16'hFF5D, 16'hFF5D, 16'hFF5D, 16'hFF5D, 16'hFF5E, 16'hFFDF, 16'hCDD8, 16'hD619, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE69A, 16'hEF1C, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCDD8, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F,
        16'hFFDF, 16'hCDD8, 16'hEF1C, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hD619, 16'hC596, 16'hFF9E, 16'hFF5D, 16'hFF5E, 16'hFF5E, 16'hEF1C, 16'hD619, 16'hDE59, 16'hDE59, 16'hBD55, 16'hB555, 16'hACD3, 16'h5A89, 16'hBD55, 16'hC5D7, 16'hDE99, 16'hD659, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hCE58, 16'hDEDA, 16'h9CD2, 16'h7B8E, 16'hD699, 16'hD658, 16'hD658, 16'hD659, 16'hD659, 16'hD659, 16'hD658, 16'hCE58, 16'hD659, 16'hE6DB, 16'hF75D, 16'hF75D, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE69A, 16'h2000, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB514, 16'h8B8E, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hEEDC, 16'hD658, 16'hD659, 16'hD659,
        16'hDE99, 16'hAD13, 16'h738D, 16'hDE99, 16'hCE58, 16'hD659, 16'hA492, 16'h9C51, 16'hD659, 16'hE69A, 16'h7B8D, 16'h9C92, 16'hEEDB, 16'hAC92, 16'hCDD7, 16'hE69A, 16'hF75D, 16'hFF5D, 16'hFF5D, 16'hFF5D, 16'hFF5D, 16'hFF9F, 16'hCDD7, 16'hDE9B, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hDE9A, 16'hEF1C, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCDD7, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD659, 16'hDE9B, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE69A, 16'hBD56, 16'hFF9E, 16'hFF5D, 16'hFF5D, 16'hFF5E, 16'hDE5A, 16'hD619, 16'hD619, 16'hE69A, 16'hC5D6, 16'h41C6, 16'h7B8E, 16'hCE18, 16'hDE59, 16'hB514, 16'hA4D2, 16'hE6DA, 16'hD659, 16'hCE58, 16'hD658, 16'hCE58, 16'hCE58, 16'hCE58, 16'hD699, 16'hBDD6, 16'h734D, 16'hCE58, 16'hD699, 16'hD658, 16'hD658, 16'hD659,
        16'hD658, 16'hCE58, 16'hD659, 16'hE6DB, 16'hF75D, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD659, 16'h2082, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC5D7, 16'h6A8A, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hF71C, 16'hD659, 16'hD658, 16'hD659, 16'hCE18, 16'h62CB, 16'hC5D6, 16'hDE99, 16'hB555, 16'h9C92, 16'hDE9A, 16'hD659, 16'hDE99, 16'hCDD7, 16'h41C6, 16'hDE19, 16'hACD3, 16'hDE18, 16'hDE5A, 16'hEEDC, 16'hFF5E, 16'hFF5D, 16'hFF5D, 16'hFF5D, 16'hFF9E, 16'hBD96, 16'hE6DC, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hDE59, 16'hEF1C, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF,
        16'hCDD7, 16'hF71D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE69A, 16'hDE5A, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hEEDC, 16'hB515, 16'hFF5E, 16'hFF5D, 16'hFF5E, 16'hEEDC, 16'hD619, 16'hDE59, 16'hE69A, 16'hB514, 16'h5249, 16'hA4D3, 16'hDE59, 16'hDE59, 16'hCE18, 16'hEF1C, 16'hD659, 16'hBD55, 16'hFF5E, 16'hD699, 16'hCE18, 16'hD658, 16'hCE58, 16'hD699, 16'hC5D6, 16'h630B, 16'hC5D7, 16'hD699, 16'hD658, 16'hD659, 16'hD659, 16'hCE58, 16'hCE58, 16'hE6DB, 16'hF75D, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hBD56, 16'h5249, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h6A08, 16'hEF1C, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'hDE9A, 16'hD618, 16'hDE9A, 16'h9450, 16'h9C92, 16'hD659, 16'h9410, 16'hD658, 16'hD658, 16'hD618, 16'hD658, 16'hE69A, 16'h9410, 16'h8BCF, 16'hB514, 16'hDE59, 16'hE65A, 16'hE69A, 16'hF75D, 16'hFF5D, 16'hFF5D, 16'hFF5D, 16'hFF9E, 16'hBD55, 16'hEEDC, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hDE59, 16'hEF1C, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hCDD8, 16'hEF1D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEEDC, 16'hD618, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF5E, 16'hF75D, 16'hFF5E, 16'hF71D, 16'hB4D4, 16'hFF5D, 16'hFF5E, 16'hFF5D, 16'hDE5A, 16'hDE59, 16'hE69A, 16'h9C52, 16'h41C7, 16'hBD95, 16'hDE99, 16'hD659, 16'hDE99, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hCDD8, 16'hDE59, 16'hFFDF,
        16'hDE9A, 16'hCE17, 16'hD699, 16'hCE58, 16'h62CB, 16'hBD95, 16'hDE99, 16'hD658, 16'hD658, 16'hCE58, 16'hCE58, 16'hDE9A, 16'hF75D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'h9451, 16'h7BCF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h7B0B, 16'hDE59, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hE6DB, 16'hDE99, 16'hBD96, 16'h6B0B, 16'hA4D2, 16'hAD13, 16'hE6DB, 16'hE6DB, 16'hE69A, 16'hD659, 16'hDE59, 16'hD618, 16'h41C7, 16'h9C92, 16'hE69A, 16'hDE59, 16'hE65A, 16'hF71C, 16'hFF5E, 16'hFF5D, 16'hFF5D, 16'hFF5E, 16'hBD15, 16'hEF1C, 16'hFF9F, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF,
        16'hD659, 16'hEEDC, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hCDD8, 16'hEF1C, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1D, 16'hC596, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hFF5D, 16'hFF5D, 16'hFF5D, 16'hFF5D, 16'hFF5D, 16'hB4D4, 16'hEEDC, 16'hFF5E, 16'hEEDC, 16'hDE59, 16'hDE59, 16'h83CF, 16'h6B0C, 16'hC596, 16'hD659, 16'hD659, 16'hEF1C, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hBD56, 16'hF71D, 16'hFF9E, 16'hE6DB, 16'hCE58, 16'h6B0C, 16'hAD54, 16'hDE99, 16'hD658, 16'hD658, 16'hCE58, 16'hD659, 16'hEF1C, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hDE9A, 16'h734D, 16'hB555, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h7B4D, 16'hBD15, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hF75D, 16'h8C11, 16'h5208, 16'hDE9A, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF71D, 16'hDE59, 16'hE69A, 16'hC596, 16'h6ACB, 16'hDE59, 16'hE69A, 16'hDE59, 16'hE69B, 16'hFF5E, 16'hFF5D, 16'hFF5D, 16'hFF5E, 16'hBD55, 16'hF71C, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hDE59, 16'hEEDC, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hCDD8, 16'hE6DC, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'hC596, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hFF5D, 16'hFF5D, 16'hFF5D, 16'hFF5D, 16'hF75D, 16'hFF5E, 16'hBD55, 16'hE6DB, 16'hFF5E, 16'hEE9B, 16'hCDD7, 16'h6ACB, 16'h7B4D,
        16'hC5D6, 16'hD659, 16'hE6DB, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'hBD55, 16'hFF9F, 16'hEF1C, 16'h630B, 16'hAD13, 16'hDE9A, 16'hCE58, 16'hD658, 16'hD658, 16'hE71B, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'hCE18, 16'h5248, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC5D7, 16'h8BCF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h3104, 16'hEF1C, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'hDE59, 16'hEE9A, 16'hB514, 16'h7B4D, 16'hDE59, 16'hE69A, 16'hDE59, 16'hF71D, 16'hFF5D,
        16'hFF5D, 16'hFF5E, 16'hBD55, 16'hF71D, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9E, 16'hFF9F, 16'hDE59, 16'hEEDB, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hCE18, 16'hDE9B, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9E, 16'hC596, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5D, 16'hFF5D, 16'hFF5D, 16'hFF5D, 16'hF75D, 16'hFF5E, 16'hD5D8, 16'hD618, 16'hF71C, 16'hACD4, 16'h49C8, 16'hA492, 16'hDE59, 16'hAC93, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD659, 16'hDE9A, 16'h6B0C, 16'hA4D3, 16'hDE99, 16'hCE58, 16'hD658, 16'hE6DA, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hDE9A,
        16'hB514, 16'h630C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h59C7, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hAD14, 16'hB555, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hC596, 16'hACD3, 16'h6B0C, 16'h62CB, 16'hDE59, 16'hE69A, 16'hE69B, 16'hFF5D, 16'hFF5D, 16'hFF5E, 16'hBD55, 16'hEEDC, 16'hFF9E, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF9F, 16'hD618, 16'hE6DB, 16'hFF9F, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hD619, 16'hDE5A, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hCD97, 16'hF71D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5D,
        16'hFF5D, 16'hFF5D, 16'hFF5D, 16'hF75D, 16'hFF5E, 16'hF6DC, 16'hB514, 16'h9410, 16'h62CB, 16'hC596, 16'hDE9A, 16'hF75D, 16'hEF1C, 16'hBD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'h628A, 16'hAD14, 16'hD659, 16'hCE58, 16'hDE9A, 16'hF71D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE6DC, 16'hD659, 16'h734D, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h7B0C, 16'hD618, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'h838F, 16'hF75E, 16'hFFDF,
        16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE69B, 16'hC597, 16'hE69B, 16'hD618, 16'h9451, 16'h734D, 16'hDE59, 16'hE69A, 16'hEF1C, 16'hFF5E, 16'hFF9E, 16'hC556, 16'hEEDB, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF9F, 16'hD618, 16'hE69B, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hDE5A, 16'hD659, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hCD97, 16'hF6DC, 16'hFF5E, 16'hFF5D, 16'hFF5D, 16'hFF5D, 16'hFF5D, 16'hFF5D, 16'hFF1D, 16'hFF5D, 16'hFF5D, 16'hC596, 16'h5208, 16'hA492, 16'hDE59, 16'hEEDC, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hCE18, 16'hDE9A, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9E, 16'h840F, 16'h9C91, 16'hD659, 16'hDE9A, 16'hF75D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9E, 16'hD659, 16'hC5D7, 16'h4A08, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD14, 16'hA493, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hBD97, 16'hB515, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9E, 16'hB515, 16'hF75E, 16'hFFDF, 16'hEF1C, 16'hE69A, 16'hACD4, 16'h5248, 16'hBD55, 16'hE69A, 16'hE69B, 16'hF75D, 16'hC556, 16'hDE19, 16'hF71D, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hD618, 16'hE69B, 16'hFF9F, 16'hFF5E, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE69A, 16'hCDD8, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F,
        16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hFF9E, 16'hD5D8, 16'hEE9B, 16'hFF5E, 16'hFF5D, 16'hFF5D, 16'hFF5D, 16'hFF1D, 16'hF71D, 16'hFF5E, 16'hF71C, 16'h9C52, 16'h734D, 16'hCDD7, 16'hEEDB, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF79E, 16'hBD56, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'h8C10, 16'h8C10, 16'hD659, 16'hE6DB, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE9B, 16'hDE99, 16'h9491, 16'h8C51, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h5A49, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9E, 16'h734D, 16'hE6DC, 16'hFFDF, 16'hFFDF, 16'hD619, 16'hD659, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'hDE5A, 16'hB514, 16'h4187, 16'h9C51, 16'hE65A, 16'hE69B, 16'hB514, 16'hDE59, 16'hE69A, 16'hEEDB, 16'hFF5D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hD618, 16'hE69A, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF5E, 16'hFF9F, 16'hE6DB, 16'hCDD7, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hDE59, 16'hE65A, 16'hFF5E, 16'hFF5D, 16'hFF5D, 16'hFF5D, 16'hFF5E, 16'hFF9E, 16'hD659, 16'h730D, 16'h940F, 16'hDE59, 16'hF75D, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hCDD7, 16'hE6DB, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'h8C11, 16'h9C92, 16'hEF1B, 16'hF75D, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF,
        16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'hD659, 16'hD699, 16'h4A08, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h5A49, 16'hD659, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE9A, 16'h83CF, 16'hFFDF, 16'hFF9E, 16'hBD96, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9E, 16'hE6DB, 16'hD618, 16'h9C51, 16'h730C, 16'hBD56, 16'hB514, 16'hDE59, 16'hE69A, 16'hE65A, 16'hE69B, 16'hF71D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hD5D8, 16'hE69A, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E,
        16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF9F, 16'hEEDC, 16'hC596, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF9F, 16'hE69B, 16'hD618, 16'hFF5E, 16'hF71D, 16'hFF5E, 16'hFF9E, 16'hE69B, 16'h9C52, 16'h730C, 16'hBD55, 16'hDE59, 16'hCDD8, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE6DC, 16'hCDD7, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF79E, 16'h734D, 16'h9C92, 16'hF75D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hD659, 16'hDEDA, 16'hA513, 16'h738E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB555, 16'h8BD0, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'hDE9A, 16'hA4D4, 16'hBD96, 16'hEEDB, 16'hDE5A, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hF71C, 16'hACD3, 16'hA492, 16'h7B4D, 16'h5208, 16'hBD55, 16'hE69A, 16'hE69A, 16'hE65A, 16'hE65A, 16'hEF1C, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hD618, 16'hE69B, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF9E, 16'hF71D, 16'hBD56, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF9E, 16'hF71C, 16'hCD97, 16'hFF5E, 16'hFF5E, 16'hF71C, 16'hACD4, 16'h6ACB, 16'h9451, 16'hE69A, 16'hF71D, 16'hFF9F, 16'hD618, 16'hEF1D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hBD96, 16'hFF5E, 16'hFFDF, 16'hEF1C, 16'h734D,
        16'hBD96, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE6DB, 16'hD659, 16'hDE9A, 16'h5A8A, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h38C2, 16'hEEDC, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE9A, 16'hD619, 16'hFF9F, 16'h838E, 16'hA4D3, 16'hF75E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE6DC, 16'hB514, 16'hE69A, 16'hD658, 16'hB514, 16'h628A, 16'h83CF, 16'hD618, 16'hE69A, 16'hE65A,
        16'hDE59, 16'hE69B, 16'hF71D, 16'hFF9E, 16'hD5D8, 16'hE69A, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF5D, 16'hBD56, 16'hFF5E, 16'hFF9E, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hD5D8, 16'hE65A, 16'hACD3, 16'h62CA, 16'h8BCF, 16'hDE9A, 16'hF75D, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hEEDC, 16'hCE18, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hEEDC, 16'hFFDF, 16'hD659, 16'h5A49, 16'hD659, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'hD658, 16'hDEDA, 16'hAD54, 16'h738E, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'h83CF, 16'hA492, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hC596, 16'hDE9B, 16'hFFDF, 16'hC597, 16'h7B8E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hBD96, 16'hF75D, 16'hFF9E, 16'hE69A, 16'hDE59, 16'hDE59, 16'hB514, 16'h7B4D, 16'hB514, 16'hE65A, 16'hE69A, 16'hDE59, 16'hDE59, 16'hEEDC, 16'hCDD7, 16'hE69B, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hBD56, 16'hF71D, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF1D, 16'hDE5A, 16'h93D0, 16'h6B0C, 16'hB555, 16'hE6DB, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hC597, 16'hF75E,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hB555, 16'h734D, 16'hEEDC, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD659, 16'hD699, 16'hDE99, 16'h630C, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h000, 16'hE69B, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'hEEDC, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD55, 16'hF75D, 16'hFFDF, 16'hFF9F, 16'h8C10, 16'hD659, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F,
        16'hFFDF, 16'hEF1C, 16'hBD56, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hF71D, 16'hE69A, 16'hE69A, 16'hD618, 16'h9410, 16'h838E, 16'hBD55, 16'hDE59, 16'hE69A, 16'hE69A, 16'hBD55, 16'hDE59, 16'hFF5D, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hC596, 16'hE69B, 16'hFF9F, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFF9E, 16'hFF1D, 16'hDE19, 16'h9C11, 16'h6ACB, 16'h9410, 16'hC596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE5A, 16'hE69B, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hE71C, 16'h8C10, 16'hACD4, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDA, 16'hD658, 16'hDEDA, 16'hAD14, 16'h8C50, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'h734D, 16'h730D, 16'hF75D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEEDC, 16'hDE9A, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hB555, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'h6B0C, 16'hF75D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hCE18, 16'hD659, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hF75D, 16'hEEDB, 16'hE69A, 16'hC596, 16'h6ACB, 16'h834E, 16'h9C51, 16'hCDD7, 16'hBD14, 16'hD5D7, 16'hEE9A, 16'hEEDB, 16'hF71C, 16'hF75D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF5E, 16'hFFDF, 16'hDE5A, 16'hDE59, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hF6DC, 16'hD618, 16'h9C51, 16'h730C, 16'h628A, 16'hACD3, 16'hE6DB, 16'hFF5D,
        16'hC597, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF71D, 16'hCDD8, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hBD96, 16'h83D0, 16'hDE9A, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hEEDB, 16'hE6DB, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE71C, 16'hD659, 16'hDE99, 16'hD659, 16'h5ACA, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h7B4D, 16'hACD3, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'hD619, 16'hFF5E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF,
        16'hEF1C, 16'hC596, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hCDD8, 16'h8BD0, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hBD55, 16'hEF1D, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hD618, 16'hACD3, 16'hD5D8, 16'h9C51, 16'h7B4D, 16'h628A, 16'h838E, 16'hC596, 16'hD618, 16'hDE19, 16'hE69A, 16'hEE9B, 16'hF71C, 16'hFF5E, 16'hFF5D, 16'hFF5D, 16'hF75D, 16'hF71D, 16'hDE9A, 16'h9C51, 16'hD619, 16'hD659, 16'hBD56, 16'hA492, 16'h8BCF, 16'h628A, 16'h6ACB, 16'h9C92, 16'hCE18, 16'hEF1C, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hBD56, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hCDD7, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hCE18, 16'h83CF, 16'hA493, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hEEDC, 16'hE659, 16'hDE59,
        16'hF71D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'hD699, 16'hD699, 16'hDEDA, 16'h9491, 16'h8C51, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h6ACB, 16'hDE59, 16'hB514, 16'hEF1D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'hD618, 16'hF71D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE9A, 16'hCDD8, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'h9C92, 16'hC5D8, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'hB514, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hCDD7, 16'hE6DC, 16'hFFDF, 16'hF75D, 16'hE6DB, 16'hD618, 16'hACD3, 16'h730C, 16'h7B4D, 16'h7B0C, 16'h7B0C, 16'h93CF, 16'h93CF, 16'h93CF, 16'h834D, 16'h7B4D, 16'h7B0C, 16'h6ACB, 16'h6A8A, 16'h838D, 16'h834D,
        16'h8BCF, 16'hA491, 16'h8BCF, 16'hCDD8, 16'hE6DB, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hC596, 16'hEEDC, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'hF75D, 16'hD69A, 16'h9411, 16'hACD4, 16'hEF1D, 16'hCDD8, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hE65A, 16'hE65A, 16'hE659, 16'hEEDC, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD699, 16'hD699, 16'hDE99, 16'hCE58, 16'h39C7, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h8C10, 16'hFFDF, 16'hA492, 16'hD659, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF71D, 16'hCE18, 16'hE6DB, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hCE18, 16'hDE5A, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF71D, 16'h628A, 16'hD65A, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hBD96, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hC556, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF75D, 16'hEEDB, 16'hE69A, 16'hBD55, 16'hC556, 16'hB515, 16'hB514, 16'hC5D7, 16'hDE59, 16'hDE5A, 16'hE69B, 16'hEEDC, 16'hF75D, 16'hFF5E, 16'hFF9F, 16'hFF9E, 16'hCDD7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hCDD8, 16'hDE9B, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hDE5A, 16'h9411, 16'h9452, 16'hE6DC, 16'hFFDF, 16'hFF9F, 16'hC596, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69B, 16'hDE59, 16'hE65A, 16'hE659, 16'hF71C, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDEDA, 16'hD659, 16'hD659, 16'hE6DA, 16'h8C50, 16'h9492, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h62CB, 16'hE6DB, 16'hEEDC, 16'hBD96, 16'hACD4, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'hCE18, 16'hDE9A, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hC5D7, 16'hE6DC, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hD619, 16'hD659, 16'h9C51, 16'hEF1C, 16'hFFDF, 16'hE6DB, 16'hD65A, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hBD55, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFF9F, 16'hFFDF, 16'hEF1C, 16'hDE5A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF75E, 16'hC596, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD659, 16'hD659, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h9C92, 16'h8C10, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hBD96, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF5E, 16'hDE59, 16'hE65A, 16'hE659, 16'hE65A, 16'hF75D, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE6DB, 16'hD699, 16'hDEDA, 16'hDE99, 16'hCE58, 16'h41C7, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC618, 16'h83CE, 16'hFF9E, 16'hBD97, 16'hFF9F, 16'h9451, 16'hEF1D, 16'hFFDF, 16'hFF9F, 16'hF75E,
        16'hD618, 16'hD618, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hBD55, 16'hEF1D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hBD56, 16'hF75E, 16'hEF1C, 16'h730C, 16'hF75E, 16'hEF1D, 16'hEEDC, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'hC597, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE6DB, 16'hCE18, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hC596, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE69B, 16'hCDD8, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h9452, 16'h7B8E, 16'hB555, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hF71D, 16'hBD96, 16'hFFDF, 16'hFF9F,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEEDC, 16'hDE19, 16'hE65A, 16'hE65A, 16'hE69B, 16'hF75E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hCE58, 16'h9451, 16'h7B8E, 16'h8C50, 16'h000, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h6B0C, 16'hDE9B, 16'hE6DB, 16'hD659, 16'hFFDF, 16'hBD97, 16'hC5D7, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hD659, 16'hCDD8, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hB515, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'hBD55, 16'hFF9E, 16'hFFDF, 16'hD659, 16'h730C, 16'hEF1C, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFF9F, 16'hFFDF, 16'hE69A, 16'hD619, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE69B, 16'hD659, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hC596, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF71D, 16'hC597, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hAD14, 16'h83CF, 16'hD659, 16'hF75D, 16'hCDD7, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1D, 16'hC597, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hDE5A, 16'hDE59, 16'hDE59, 16'hE65A, 16'hEEDC, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hCE18,
        16'h6ACB, 16'h9C91, 16'hB554, 16'hD699, 16'hAD54, 16'h4A49, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hD69A, 16'h8BCF, 16'hFFDF, 16'hBD96, 16'hEF1D, 16'hFFDF, 16'hEF1C, 16'h8C10, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hD659, 16'hCDD7, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'hB515, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'hC596, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE5A, 16'h628A, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE59, 16'hE69B, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hDE9A, 16'hD659, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hC596, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hCDD8, 16'hFFDF, 16'hFF9F, 16'hBD96, 16'h734D, 16'hB555, 16'hFF9F,
        16'hFFDF, 16'hEF1C, 16'hC597, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'hC597, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'hD618, 16'hDE59, 16'hDE59, 16'hE69A, 16'hF71D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF79E, 16'hA493, 16'h9C52, 16'hEEDC, 16'hE6DA, 16'hA4D2, 16'hD699, 16'hDEDA, 16'h5289, 16'hC5D7, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h734D, 16'hDE9A, 16'hF75D, 16'hBD96, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'h9C51, 16'hDE9A, 16'hFFDF, 16'hFF9F, 16'hDE9A, 16'hC596, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'hBD56, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE69B, 16'hCDD8,
        16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'h7B8E, 16'hB555, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD618, 16'hEF1D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD65A, 16'hDE9A, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hBD96, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9E, 16'hCE18, 16'h7B8E, 16'hACD4, 16'hEF1D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE6DB, 16'hCDD8, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE6DC, 16'hC597, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEEDC, 16'hD618, 16'hDE59, 16'hDE59, 16'hEEDB, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hDEDB, 16'h8BCF, 16'hCE19, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'hA512, 16'hB595, 16'hE71B, 16'hB555, 16'h630C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h730C, 16'hFFDF, 16'hCE18, 16'hD659, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hCE18, 16'hB515, 16'hFFDF, 16'hFFDF, 16'hDE9B, 16'hBD55, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE6DB, 16'hCDD7, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE5A, 16'hD659, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hB555, 16'h734D, 16'hE6DC, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hD618, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD659, 16'hE6DB, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hBD96, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hD659, 16'h9451, 16'hAD14, 16'hE6DC, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE69B, 16'hD619, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE6DB, 16'hC597, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'hD618, 16'hDE19, 16'hE69A, 16'hF71C, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hC5D7, 16'h9411, 16'hEF1C, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hBDD6, 16'h94D2, 16'hDEDA, 16'hD659, 16'h4A48, 16'hD69A, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h738E, 16'hCE18, 16'hFFDF, 16'hB555, 16'hF75D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'h9410, 16'hF75E, 16'hFFDF, 16'hE6DB, 16'hB514, 16'hF75D, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE5A, 16'hCE18, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hCDD8, 16'hDE9A, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hDE9A, 16'h83CF, 16'hAD15, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hE69B, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD659, 16'hE6DC, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC596, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9B, 16'h9451, 16'h9451, 16'hDE9B, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE9A, 16'hD659, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE69B, 16'hC597, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hD618, 16'hD618,
        16'hD619, 16'hEF1C, 16'hFF5D, 16'hFF5E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'hA493, 16'hC596, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hDE99, 16'h8450, 16'hCE58, 16'hE6DB, 16'hA4D3, 16'h8410, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD69A, 16'h6B0C, 16'hFFDF, 16'hE6DC, 16'hB555, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hB515, 16'hCDD8, 16'hFFDF, 16'hEF1C, 16'hAD14, 16'hF71D, 16'hFF5E, 16'hFF9E, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD619, 16'hD659, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hC596, 16'hEEDC, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hB515, 16'h8BCF, 16'hD619, 16'hFF9F, 16'hFFDF, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD619, 16'hEEDC, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hCDD7, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD65A, 16'h8C10, 16'h8BCF, 16'hBD96, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD619, 16'hDE5A, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE9B, 16'hCDD7, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'hD5D8, 16'hDE19, 16'hE69A, 16'hF75D, 16'hF75D, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE6DB, 16'h9410, 16'hDE9B, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hEF1B, 16'h9D12, 16'hBDD6, 16'hDEDA, 16'hD658, 16'h39C6, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h7B8E, 16'hBD96, 16'hFFDF, 16'hD659, 16'hCE18, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'h9C51, 16'hFFDF, 16'hF75D, 16'hACD3, 16'hEF1C, 16'hF75D, 16'hF75D, 16'hFF5E, 16'hFF9F, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hC5D7, 16'hDE9B, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD55, 16'hF75D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hEF1D, 16'hA492, 16'h8BD0, 16'hDE5A, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD619, 16'hEEDC, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD659, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hCE19, 16'h7B8E, 16'h83CF, 16'hE6DB, 16'hEF1C, 16'hD619, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD619, 16'hDE9B, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE9A, 16'hCE18, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE6DB, 16'hCDD8, 16'hD619, 16'hEF1C, 16'hFF5D, 16'hFF5D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hD659, 16'h7B4D, 16'hEF1D, 16'hFFDF, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'hB595, 16'hA554, 16'hDE9A, 16'hDEDA, 16'h7B8E, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9B, 16'h5A8A, 16'hFF9E, 16'hFFDF, 16'hBD96, 16'hE6DC, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hACD4, 16'hE69B, 16'hF75E, 16'hACD3, 16'hEEDB, 16'hEF1C, 16'hF75D, 16'hF75D, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hBD96, 16'hE6DC, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hB514, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hE69B, 16'h9C51, 16'h93D0, 16'hCDD8, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hD659, 16'hEEDB, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hF75D, 16'hCE18, 16'h83CF, 16'h9C92, 16'hDE9A, 16'hFF9F, 16'hFFDF, 16'hDE9B, 16'hCE18, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hCDD8, 16'hE6DB, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD659, 16'hCE18, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hDE59, 16'hCDD7, 16'hE69B, 16'hFF5D, 16'hF75D, 16'hFF5E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hC5D8, 16'h7B8E, 16'hF75E, 16'hFFDF, 16'hFF9E, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF75E, 16'hCE17, 16'h9D13, 16'hD699, 16'hDE9A, 16'hC617,
        16'h4A48, 16'hF79D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9451, 16'hB555, 16'hFFDF, 16'hFF9E, 16'hB555, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hEF1C,
        16'hEF1C, 16'hFFDF, 16'hDE9A, 16'hB514, 16'hF75E, 16'hAD13, 16'hEEDB, 16'hEF1C, 16'hEF1C, 16'hF71D, 16'hF75D, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hB555, 16'hEF5D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hB555, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE9A, 16'hD619, 16'hC597, 16'h7B4D, 16'h9C52, 16'hCE18, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE9A, 16'hE6DB, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1D, 16'hB556, 16'h8C10, 16'hA4D4, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE5A, 16'hD659, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hC5D7, 16'hE6DC, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF,
        16'hD659, 16'hD659, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hCDD8, 16'hD618, 16'hF71D, 16'hFF5D, 16'hF75D, 16'hFF5E, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hB555, 16'h83CF, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE9A, 16'hF75D, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hDE99, 16'hA513, 16'hC617, 16'hD699, 16'hDEDA, 16'h734D, 16'hB596, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE6DB, 16'h5A48, 16'hF71D, 16'hFFDF, 16'hE6DC, 16'hBD56, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hCE18, 16'hE6DC, 16'hFFDF, 16'hFF9E, 16'hACD4, 16'hE6DB, 16'hAD14, 16'hE6DB, 16'hEF1C, 16'hEEDC, 16'hEEDC, 16'hEF1C, 16'hF75D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hB515, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hEF1D, 16'hBD56, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC597, 16'hEF1D, 16'hFFDF, 16'hF75E, 16'hCE19, 16'hA4D3, 16'h8BCF, 16'h9C51, 16'hC5D7, 16'hE6DB, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFF5E, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hD65A, 16'hA493, 16'h8BCF, 16'hBD96, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hD618, 16'hD65A, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hC596, 16'hEF1C, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD619, 16'hD65A, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hF75D, 16'hC596, 16'hE69B, 16'hFF5D, 16'hF75D, 16'hF75D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hB555, 16'h9451, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hEF1C,
        16'hDE9B, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE6DB, 16'hBDD6, 16'hCE58, 16'hDEDA, 16'hE6DA, 16'hC5D7, 16'h630C, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'h9451, 16'h9C51, 16'hFFDF, 16'hFFDF, 16'hD619, 16'hCE19, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hC597, 16'hF75E, 16'hFF9F, 16'hFFDF, 16'hCE19, 16'hBD96, 16'hB555, 16'hE6DB, 16'hEF1C, 16'hEF1C, 16'hEEDC, 16'hEF1C, 16'hEF1C, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hAD14, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE6DC, 16'hC597, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hB555, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'hDE9A, 16'hCDD8, 16'h9C51, 16'h8C10, 16'h9410, 16'hB514, 16'hBD56, 16'hCDD8, 16'hDE9A, 16'hD65A, 16'hD65A, 16'hCE18, 16'hBD56, 16'h9C51, 16'h7B8E, 16'hA492, 16'hD659, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hC5D7, 16'hDE9B, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD56, 16'hEF1D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hCDD8, 16'hDE5A, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hEEDB, 16'hC596, 16'hF71D, 16'hF75D, 16'hF75D, 16'hF75D, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hB515, 16'h9411, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hCE18, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'hDE99, 16'hBDD6, 16'hA513, 16'hB554, 16'hA4D2, 16'h000, 16'hD659, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h51C7, 16'hE6DB, 16'hFFDF, 16'hFFDF, 16'hC597, 16'hE6DB, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'hC597, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'h9C92, 16'hB514, 16'hE6DB, 16'hEF1C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEF1C, 16'hEF1D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'hB555, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F,
        16'hFFDF, 16'hDE9A, 16'hCDD8, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hBD55, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hD619, 16'hF75D, 16'hE6DC, 16'hD659, 16'hBD96, 16'h9C93, 16'h9C92, 16'h9451, 16'h9C92, 16'hA4D3, 16'hAD15, 16'hD659, 16'hF75E, 16'hFFDF, 16'hF75D, 16'hCE18, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hC5D7, 16'hE6DC, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hB515, 16'hF75D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hC597, 16'hDE9B, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9F, 16'hDE59, 16'hD618, 16'hF75D, 16'hF75D, 16'hF75D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F,
        16'hFF9F, 16'hFFDF, 16'hB555, 16'h8C10, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD659, 16'hEF1C, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hDE9A, 16'h840F, 16'h6B4C, 16'h7BCE, 16'hBD95, 16'hBDD6, 16'h840F, 16'h8C50, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9C92, 16'h8BCF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hBD56, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE69B, 16'hCDD8, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hBD56, 16'h9C51, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'hBD55, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD619, 16'hD659, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1D, 16'hB555, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hBD56, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hDE9B, 16'hCE18, 16'hFFDF, 16'hFF9F,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hC596, 16'hEF1C, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hB515, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hBD96, 16'hE6DB, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hCDD7, 16'hE69B, 16'hF75D, 16'hF75D, 16'hFF5D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hC5D8, 16'h8C10, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'hE69B, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9E, 16'h9C93, 16'h8BD0, 16'hB555, 16'hD658, 16'hA4D2, 16'hCE58, 16'hDEDA, 16'hCE58, 16'h41C7, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h000, 16'hCDD7, 16'hFF9F, 16'hFF9F, 16'hF75D, 16'hBD56, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hD659, 16'hDE5A, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE6DB, 16'h83CF, 16'hEEDB, 16'hEF1C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEF1D, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE6DB, 16'hBD96, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hCDD8, 16'hE69B, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEEDC, 16'hBD96, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'hBD56, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hDE9A, 16'hCE18, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hBD96, 16'hEF5D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hB515, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hC596, 16'hEEDC, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E,
        16'hC596, 16'hEEDC, 16'hF75D, 16'hF75D, 16'hFF5E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hCE59, 16'h7B4D, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hE6DC, 16'h83D0, 16'hBD97, 16'hFF9F, 16'hFF9E, 16'hE6DA, 16'h9CD2, 16'hBDD6, 16'hD699, 16'hDEDA, 16'h7BCF, 16'hA514, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'h9C92, 16'h2800, 16'hF6DC, 16'hFF9E, 16'hFFDF, 16'hE69B, 16'hC5D7, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hC597, 16'hE6DB, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hA4D3, 16'hE69A, 16'hEF1C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEF1C, 16'hEF1C, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE9A, 16'hC5D7, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hBD96, 16'hE6DC, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hE69B, 16'hC597, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF71D, 16'hBD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD659, 16'hD619, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD55, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hB515, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hBD55, 16'hEF1D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hF71C, 16'hBD55, 16'hF71D, 16'hF75D, 16'hF75D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'h730C, 16'hEF1C, 16'hEEDC, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hEF1D, 16'hC5D8, 16'hB555, 16'hDE9B, 16'hFFDF, 16'hFF9F, 16'hFF9E, 16'hE6DB, 16'hAD13, 16'hAD54, 16'hDE9A, 16'hDE9A, 16'hAD54, 16'h39C7, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h6A8A, 16'h93CF, 16'hF71D, 16'hFF5E, 16'hFF9F, 16'hD659, 16'hDE5A, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hBD96, 16'hF75D, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hC596, 16'hDE5A, 16'hEF1C,
        16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEF1C, 16'hEF1C, 16'hF75D, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD619, 16'hCE18, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hBD55, 16'hEF1D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD659, 16'hCE18, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1D, 16'hC5D7, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hCDD8, 16'hDE5A, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hBD56, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'hB555, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB555, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hDE9A, 16'hBD56, 16'hFF5E, 16'hF75D, 16'hF75D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'h6B0C, 16'hE6DB, 16'hFFDF, 16'hDE59, 16'hF75D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hC5D8, 16'hBD56, 16'h838E, 16'hEF1D, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hEF1C, 16'hB595, 16'h9CD2, 16'hDE9A, 16'hDE99, 16'hC617, 16'h000, 16'hCE59, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA4D3, 16'hAC93, 16'h9C11, 16'hEEDC, 16'hFF9E, 16'hFF9F, 16'hC596, 16'hEEDC, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hBD55, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9F, 16'hAD14, 16'hD659, 16'hEF1C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEF1C, 16'hEF1C, 16'hEF1C, 16'hF71D, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hC5D7, 16'hD619, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hBD55, 16'hF75D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD619, 16'hDE5A, 16'hFFDF, 16'hFF9F,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'hCDD7, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hC596, 16'hDE9B, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9E, 16'hBD56, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF71D, 16'hB555, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hBD55, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hF75D, 16'hFF9E, 16'hCDD8, 16'hCDD8, 16'hFF5E, 16'hF75D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'h838E, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hEF1D, 16'hCE18, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9E, 16'hA493, 16'hB555, 16'hFFDF, 16'hC5D8, 16'hCE18, 16'hFFDF, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hF75D, 16'hC5D6, 16'h8C50, 16'hD699, 16'hD699, 16'hD699, 16'h4A48, 16'h738D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF1C, 16'h7B0C, 16'hFF5E, 16'hA492, 16'hDE5A, 16'hFF9F, 16'hFF5E, 16'hBD56, 16'hF75D, 16'hFFDF, 16'hFF9F,
        16'hFFDF, 16'hF75D, 16'hC596, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hA4D3, 16'hD618, 16'hEF1C, 16'hEEDC, 16'hEEDC, 16'hEEDC, 16'hEF1C, 16'hEF1C, 16'hEF1C, 16'hEF1C, 16'hFF9E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hBD96, 16'hDE9A, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hAD14, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hC5D7, 16'hE69B, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE6DB, 16'hCE18, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hBD96, 16'hE6DC, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'hBD56, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'hB555, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hBD55, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hF75D, 16'hFF5E, 16'hB514, 16'hDE59, 16'hFF5E, 16'hF75D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hA4D3, 16'hC597, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hC5D7, 16'hEF1D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'h83CF, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hE69B, 16'hB555, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF75E, 16'hCE18, 16'h8C10, 16'hD659, 16'hD699, 16'hDE99, 16'h8410, 16'h000, 16'hDEDB, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hA4D3, 16'hB515, 16'hFFDF, 16'hC597, 16'hACD3, 16'hFFDF, 16'hF71D, 16'hC556, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE6DC, 16'hC5D7, 16'hFFDF, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hA493, 16'hCE18, 16'hEF1C, 16'hEEDC, 16'hEF1C, 16'hEF1C, 16'hEF1C, 16'hEF1C, 16'hF71D, 16'hF71D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hBD56, 16'hE6DB, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hAD14, 16'hFF9E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hC596, 16'hEF1C, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE9A, 16'hD618, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hBD55, 16'hEF1D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1D, 16'hBD96, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEEDC, 16'hBD56, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'hB555, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hF75E, 16'hF75D, 16'hFF5D, 16'hF75D, 16'hF71D, 16'hA492, 16'hEEDB, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hC597, 16'hA4D4, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE6DB, 16'hCE18, 16'hFFDF, 16'hFF9F, 16'hFF9F,
        16'hFFDF, 16'hD659, 16'h7B8E, 16'hE6DB, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'hAD14, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hD659, 16'h8C50, 16'hC617, 16'hD699, 16'hDE99, 16'hAD14, 16'h734D, 16'h8C51, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hEF5D, 16'h730C, 16'hF75D, 16'hFF9F, 16'hF75D, 16'h8BCF, 16'hF71D, 16'hF71C, 16'hCDD8, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFFDF, 16'hDE9B, 16'hD618, 16'hFFDF, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF9F, 16'h9C92, 16'hCDD7, 16'hEF1C, 16'hEEDB, 16'hEF1C, 16'hEF1C, 16'hF71C, 16'hF71C, 16'hF71D, 16'hF71D, 16'hF75D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hB555, 16'hEF1C, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF71D, 16'hAD14, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hBD96, 16'hF71D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD65A, 16'hD619, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB515, 16'hF75D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'hC5D7, 16'hFFDF,
        16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE6DC, 16'hBD96, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'hBD55, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hF75E, 16'hF75D, 16'hF75D, 16'hFF5E, 16'hEEDC, 16'h9C11, 16'hF71C, 16'hFF5D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE6DB, 16'h72CB, 16'hE69B, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hBD96, 16'hEF1D, 16'hFFDF, 16'hFFDF, 16'hBD96, 16'h83CF, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD14, 16'hF75D, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hE6DB, 16'h9491, 16'hBDD6, 16'hDE9A, 16'hDE9A, 16'hB595, 16'hAD14, 16'h5ACB, 16'hE71C, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD14, 16'hB515, 16'hFFDF, 16'hFF9E, 16'hFFDF, 16'hCDD8, 16'hBD96, 16'hEEDC, 16'hD619, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFFDF, 16'hD659, 16'hDE9A, 16'hFFDF, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'h9451, 16'hC5D7, 16'hEF1C, 16'hEEDB, 16'hEF1C, 16'hEF1C, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF75D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hAD14, 16'hEF1D,
        16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hEEDC, 16'hAD14, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hBD56, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD659, 16'hDE5A, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hB514, 16'hF75E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE6DB, 16'hC5D7, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE9B, 16'hC596, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1D, 16'hBD56, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hF75E, 16'hF75D, 16'hF75D, 16'hF75D, 16'hFF5E, 16'hD619, 16'hA492, 16'hFF5E, 16'hF75D, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'h7B8E,
        16'hEEDC, 16'hD659, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEEDC, 16'hEF1C, 16'hFFDF, 16'hAD14, 16'h9C92, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hB555, 16'hE6DC, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hEF1C, 16'hA513, 16'hB595, 16'hDE9A, 16'hDE9A, 16'hBDD6, 16'hB595, 16'h9492, 16'h9CD3, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hEF5D, 16'h628A, 16'hEF1D, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hB515, 16'hC596, 16'hEF1C, 16'hFF9F, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hCDD8, 16'hE6DB, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF9F, 16'h9451, 16'hC5D7, 16'hEF1C, 16'hEEDC, 16'hEF1C, 16'hF71C, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF75D, 16'hF75D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hB514, 16'hF75E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE6DC, 16'hB555, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hB515, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD619, 16'hDE9A, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9E,
        16'hB514, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE9B, 16'hC5D7, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE9A, 16'hC5D7, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE6DC, 16'hC596, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hF75E, 16'hF75D, 16'hF75D, 16'hF71D, 16'hFF9E, 16'hC596, 16'hB514, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'h8C10, 16'hC5D8, 16'hFFDF, 16'hCE18, 16'hEF1C, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF5E, 16'h9C52, 16'hB556, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hC597, 16'hDE5A, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hEF1C, 16'hB555, 16'hA514, 16'hDE9A, 16'hD699, 16'hC617, 16'hAD54, 16'hCE58, 16'h4208, 16'hEF5D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hAD14, 16'hA4D3, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hF75E, 16'hACD3, 16'h838E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hC5D7, 16'hF71D, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'h9410, 16'hC596, 16'hEF1C, 16'hEEDC, 16'hF71C, 16'hF71D, 16'hF71D, 16'hF71D, 16'hF75D, 16'hF75D, 16'hF75D,
        16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFF5E, 16'hAD14, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hDE9B, 16'hBD96, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF75E, 16'hB515, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hCDD8, 16'hE69A, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'hB515, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE9A, 16'hCE19, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE5A, 16'hCDD8, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE69B, 16'hC5D7, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hF75D, 16'hF75D,
        16'hF75D, 16'hFF9E, 16'hA4D3, 16'hC596, 16'hFF9E, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hC5D7, 16'h9451, 16'hFFDF, 16'hFFDF, 16'hE6DC, 16'hCE18, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hDE9A, 16'hA493, 16'hD65A, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD619, 16'hCDD8, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF75D, 16'hC5D6, 16'h9CD2, 16'hDE9A, 16'hD699, 16'hD699, 16'hA4D3, 16'hDE9A, 16'h83CF, 16'hAD54, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hF75E, 16'h6A8B, 16'hEF1D, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hC5D7, 16'hE6DB, 16'h9451, 16'hF71D, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hC596, 16'hFF5E, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'h9C91, 16'hB555, 16'hEF1C, 16'hEF1C, 16'hF71D, 16'hF71D, 16'hF75D, 16'hF75D, 16'hF75D, 16'hF75D, 16'hF75D, 16'hF75D, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hF75D, 16'hB515, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hDE5A, 16'hC596, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF75D, 16'hBD55, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hCDD7, 16'hE6DB, 16'hFFDF,
        16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1D, 16'hBD96, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE5A, 16'hD659, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD659, 16'hCE18, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE9A, 16'hCDD8, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hF75D, 16'hF75D, 16'hF75D, 16'hFF5E, 16'h9411, 16'hD618, 16'hFF9E, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hE6DC, 16'h8C10, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hCDD8, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hD659, 16'h72CC, 16'hE6DB, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE9B, 16'hC597, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hCE58, 16'h9451, 16'hD659, 16'hD699, 16'hDEDA,
        16'hA513, 16'hC5D7, 16'hCE18, 16'h4207, 16'hF75D, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hB555, 16'h9411, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hF71D, 16'hCE18, 16'hFFDF, 16'hAD14, 16'hCDD8, 16'hFFDF, 16'hFF9E, 16'hFF9F, 16'hF75D, 16'hCD97, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E,
        16'hFF9E, 16'h9C51, 16'hBD55, 16'hEF1C, 16'hEF1C, 16'hF71D, 16'hF71D, 16'hF75D, 16'hF75D, 16'hF75D, 16'hF75D, 16'hF75D, 16'hFF5D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hEF1D, 16'hB515, 16'hFF9F, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hD619, 16'hC597, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hEF1D, 16'hBD56, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hC597, 16'hE6DB, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE6DC, 16'hBD96, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD659, 16'hDE5A, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hD619, 16'hD618, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE9A, 16'hCE18, 16'hFFDF, 16'hFF9F, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hF75D, 16'hFF5D, 16'hF71D, 16'h8B8F, 16'hE69B, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'h9411, 16'hDE9B, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE6DC, 16'hF71D, 16'hFFDF, 16'hFFDF, 16'hCE18, 16'h8BD0, 16'hEF1D, 16'hDE5A, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'hB555, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hDE9A, 16'h8C50, 16'hCE58, 16'hD699, 16'hDE9A, 16'hB555, 16'hAD13, 16'hE6DB, 16'h7B8E, 16'hB595, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'h6ACB, 16'hDE9B, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hEEDC, 16'hEEDC, 16'hFFDF, 16'hDE5A, 16'h8C10, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hF71D, 16'hCDD7, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hA4D2, 16'hB555, 16'hEEDC, 16'hEF1C, 16'hF75D, 16'hF71D, 16'hF75D, 16'hF75D, 16'hF75D, 16'hF75D, 16'hFF5D, 16'hFF5D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hEEDC, 16'hB555, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hD619, 16'hCDD8, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE6DC,
        16'hC596, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hBD56, 16'hEF1C, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hE69B, 16'hC5D7, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hD618, 16'hDE9A, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hD619, 16'hD619, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hD659, 16'hD618, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hF75D, 16'hFF5E, 16'hE6DB, 16'h8BCF, 16'hF71D, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hBD96, 16'hB514, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hBD96, 16'h9C92, 16'hF75E, 16'hFFDF, 16'hBD96, 16'hF75E, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF,
        16'hF75E, 16'hACD4, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hE6DB, 16'h9491, 16'hC617, 16'hDE9A, 16'hDE9A, 16'hC5D7, 16'h9491, 16'hE6DB, 16'hC617, 16'h4208, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD97, 16'h83CF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hDE9A, 16'hF71D, 16'hFFDF, 16'hFF5E,
        16'h838F, 16'hEF1D, 16'hFF9F, 16'hFFDF, 16'hEEDC, 16'hD5D8, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hAD13, 16'hAD14, 16'hEEDB, 16'hEF1C, 16'hF75D, 16'hF75D, 16'hF75D, 16'hF75D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5D, 16'hFF5E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hEF1C, 16'hC5D7, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hCDD8, 16'hCDD8, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE69B, 16'hCDD8, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hBD55, 16'hEF1D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hDE9A, 16'hCE18, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hCDD7, 16'hDE9B, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF,
        16'hD619, 16'hDE5A, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hD619, 16'hD65A, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hF75D, 16'hFF9E, 16'hD659, 16'h9450, 16'hFF9E, 16'hFF9F, 16'hFFDF, 16'hE6DC, 16'h8C10, 16'hE6DC, 16'hE6DB, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hAD14, 16'hBD56, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hC5D8, 16'hDE9B, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hB515, 16'hF79E, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hEF1C, 16'h9CD2, 16'hBD96, 16'hDEDA, 16'hD699, 16'hCE58, 16'h8C50, 16'hD699, 16'hDEDA, 16'h6B4D, 16'hAD55, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF,
        16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'h730C, 16'hD65A, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hC597, 16'hF71D, 16'hFF9F, 16'hFFDF, 16'hACD3, 16'hC5D8, 16'hFFDF, 16'hFFDF, 16'hE69B, 16'hD619, 16'hFF9F, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9F, 16'hB514, 16'hACD3, 16'hEEDC, 16'hEF1C, 16'hF75D, 16'hF75D, 16'hF75D, 16'hF75D, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF9E, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hE6DC, 16'hC5D7, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hCDD7, 16'hCE18, 16'hFFDF, 16'hFF9F,
        16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hDE9B, 16'hCE18, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hB514, 16'hF75D, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hD659, 16'hD659, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hC5D7, 16'hE6DB, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hD659, 16'hD659, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hCDD8, 16'hDE9A, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hFF9E, 16'hFF9E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hFF5E, 16'hF75D, 16'hFF9E, 16'hC597, 16'hACD3, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'h9411, 16'hDE9A, 16'hFFDF, 16'hCE18, 16'hFFDF, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFFDF, 16'hBD55, 16'hC5D7, 16'hFFDF, 16'hFF9F, 16'hFF9F,
        16'hFFDF, 16'hDE9A, 16'hCE18, 16'hFFDF, 16'hFF9F, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hBD96, 16'hF75D, 16'hFFDF, 16'hFF9F, 16'hFF9F, 16'hFF9F, 16'hF75D, 16'hAD14, 16'hB555, 16'hDEDA, 16'hD699, 16'hD699, 16'h9451, 16'hCE58, 16'hE6DA, 16'hBDD6, 16'h5A8A, 16'hF79E, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF, 16'hFFDF
    };
endmodule

/****************************************************************************************************************/
module m_st7789_display(w_clk, st7789_SDA, st7789_SCL, st7789_DC, st7789_RES, w_raddr, w_rdata, w_mode);
    input  wire w_clk; // main clock signal (100MHz)
    output wire st7789_SCL;
    inout  wire st7789_SDA;
    output wire st7789_DC;
    output wire st7789_RES;
    output wire [15:0] w_raddr;
    input  wire [15:0] w_rdata;
    input  wire [1:0] w_mode;

    wire w_clk_t = w_clk;

    reg [31:0] r_cnt=1;
    always @(posedge w_clk_t) r_cnt <= (r_cnt==0) ? 0 : r_cnt + 1;
    reg r_RES = 1;
    always @(posedge w_clk_t) begin
        if      (r_cnt==10_000) r_RES <= 0;
        else if (r_cnt==20_000) r_RES <= 1;
    end
    assign st7789_RES = r_RES;

    wire busy;
    reg r_en = 0;
    reg init_done = 0;
    reg [4:0]  r_state  = 0;
    reg [19:0] r_state2 = 0;

    reg [8:0] r_dat = 0;

    reg [15:0] r_c = 16'hf800;
    reg [15:0] r_pagecnt = 0;

    always @(posedge w_clk_t) if(!init_done) begin
        r_en <= (r_cnt>30_000 && !busy && r_cnt[10:0]==0);
    end else begin
        r_en <= (!busy);
    end

    always @(posedge w_clk_t) if(r_en && !init_done) r_state  <= r_state  + 1;

    always @(posedge w_clk_t) if(r_en &&  init_done) begin
        r_state2 <= (r_state2==115210) ? 0 : r_state2 + 1; // 11 + 240x240*2 = 11 + 115200 = 115211
        if(r_state2==115210) r_pagecnt <= r_pagecnt + 1;
    end

    reg [7:0] r_x = 0;
    reg [7:0] r_y = 0;
    always @(posedge w_clk_t) if(r_en &&  init_done && r_state2[0]==1) begin
       r_x <= (r_state2<=10 || r_x==239) ? 0 : r_x + 1;
       r_y <= (r_state2<=10) ? 0 : (r_x==239) ? r_y + 1 : r_y;
    end

    wire [7:0] w_nx = 239-r_x;
    wire [7:0] w_ny = 239-r_y;
    assign w_raddr = (w_mode==0) ? {r_y, r_x} :  // default
                     (w_mode==1) ? {r_x, w_ny} : // 90 degree rotation
                     (w_mode==2) ? {w_ny, w_nx} : {w_nx, r_y} ; //180 degree, 240 degree rotation

    reg  [15:0] r_color = 0;
    always @(posedge w_clk_t) r_color <= w_rdata;

    always @(posedge w_clk_t) begin
        case (r_state2) /////
            0:  r_dat<={1'b0, 8'h2A};     //
            1:  r_dat<={1'b1, 8'h00};     //
            2:  r_dat<={1'b1, 8'h00};     //
            3:  r_dat<={1'b1, 8'h00};     //
            4:  r_dat<={1'b1, 8'd239};    //
            5:  r_dat<={1'b0, 8'h2B};     //
            6:  r_dat<={1'b1, 8'h00};     //
            7:  r_dat<={1'b1, 8'h00};     //
            8:  r_dat<={1'b1, 8'h00};     //
            9:  r_dat<={1'b1, 8'd239};    //
            10: r_dat<={1'b0, 8'h2C};     //
            default: r_dat <= (r_state2[0]) ? {1'b1, r_color[15:8]} :{ 1'b1, r_color[7:0]};
        endcase
    end

    reg [8:0] r_init = 0;
    always @(posedge w_clk_t) begin
        case (r_state) /////
            0:  r_init<={1'b0, 8'h01};  //
            1:  r_init<={1'b0, 8'h11};  //
            2:  r_init<={1'b0, 8'h3A};  //
            3:  r_init<={1'b1, 8'h55};  //
            4:  r_init<={1'b0, 8'h36};  //
            5:  r_init<={1'b1, 8'h00};  //
            6:  r_init<={1'b0, 8'h2A};  //
            7:  r_init<={1'b1, 8'h00};  //
            8:  r_init<={1'b1, 8'h00};  //
            9:  r_init<={1'b1, 8'h00};  //
            10: r_init<={1'b1, 8'd240}; //
            11: r_init<={1'b0, 8'h2B};  //
            12: r_init<={1'b1, 8'h00};  //
            13: r_init<={1'b1, 8'h00};  //
            14: r_init<={1'b1, 8'h00};  //
            15: r_init<={1'b1, 8'd240}; //
            16: r_init<={1'b0, 8'h21};  //
            17: r_init<={1'b0, 8'h13};  //
            18: r_init<={1'b0, 8'h29};  //
            19: init_done <= 1;
        endcase
    end

    wire [8:0] w_data = (init_done) ? r_dat : r_init;
    m_spi spi0 (w_clk_t, r_en, w_data, st7789_SDA, st7789_SCL, st7789_DC, busy);
endmodule


/****** SPI send module,  SPI_MODE_2, MSBFIRST                                        *****/
/******************************************************************************************/
module m_spi(w_clk, en, d_in, SDA, SCL, DC,  busy);
    input  wire w_clk;       // 100KHz input clock !!
    input  wire en;          // enable
    inout  wire SDA;         //
    output wire SCL;         //
    output wire DC;          //
    input  wire [8:0] d_in;  // 1-bit data/control & 8-bit data
    output wire busy;        // busy

    reg [5:0] r_state=0;  //
    reg [7:0] r_cnt=0;    //
    reg r_SCL = 1;        //
    reg r_SDA = 1;        //
    reg r_DC  = 0;        // Data/Control
    reg [7:0] r_data = 0; //

    always @(posedge w_clk) begin
        if(en && r_state==0) begin
            r_state <= 1;
            r_data  <= d_in[7:0];
            r_DC    <= d_in[8];
            r_SDA   <= 0;
            r_cnt   <= 0;
        end
        else begin
            r_cnt <= (r_state==0) ? 0 : r_cnt + 1;
            if(r_state!=0 && r_cnt==18) r_state <= 0;
            if(r_cnt>0 && r_cnt[0]==0) r_data <= {r_data[6:0], 1'b0};
        end
    end

    always @(posedge w_clk) if(r_state!=0 && (r_cnt>=1) && (r_cnt<=16)) r_SCL <= ~r_SCL;

    assign SDA = r_data[7];
    assign SCL = r_SCL;
    assign DC  = r_DC;
    assign busy = (r_state!=0 || en);
endmodule
/******************************************************************************************/